MACRO DP_NMOS_B_83449181_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_83449181_X1_Y1 0 0 ;
  SIZE 5160 BY 9240 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 7420 3180 7700 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 1120 2320 1400 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 1540 3180 1820 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 5320 2320 5600 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 5740 3180 6020 ;
    END
  END GB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1550 1960 3610 2240 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 2025 1175 2275 4705 ;
    LAYER M1 ;
      RECT 2025 4955 2275 5965 ;
    LAYER M1 ;
      RECT 2025 7055 2275 8065 ;
    LAYER M1 ;
      RECT 1595 1175 1845 4705 ;
    LAYER M1 ;
      RECT 2455 1175 2705 4705 ;
    LAYER M1 ;
      RECT 2885 1175 3135 4705 ;
    LAYER M1 ;
      RECT 2885 4955 3135 5965 ;
    LAYER M1 ;
      RECT 2885 7055 3135 8065 ;
    LAYER M1 ;
      RECT 3315 1175 3565 4705 ;
    LAYER V1 ;
      RECT 2065 1175 2235 1345 ;
    LAYER V1 ;
      RECT 2065 5375 2235 5545 ;
    LAYER V1 ;
      RECT 2065 7475 2235 7645 ;
    LAYER V1 ;
      RECT 2925 1595 3095 1765 ;
    LAYER V1 ;
      RECT 2925 5795 3095 5965 ;
    LAYER V1 ;
      RECT 2925 7475 3095 7645 ;
    LAYER V1 ;
      RECT 1635 2015 1805 2185 ;
    LAYER V1 ;
      RECT 2495 2015 2665 2185 ;
    LAYER V1 ;
      RECT 3355 2015 3525 2185 ;
    LAYER V0 ;
      RECT 2065 3335 2235 3505 ;
    LAYER V0 ;
      RECT 2065 3675 2235 3845 ;
    LAYER V0 ;
      RECT 2065 5375 2235 5545 ;
    LAYER V0 ;
      RECT 2065 7475 2235 7645 ;
    LAYER V0 ;
      RECT 1635 3335 1805 3505 ;
    LAYER V0 ;
      RECT 1635 3675 1805 3845 ;
    LAYER V0 ;
      RECT 2495 3335 2665 3505 ;
    LAYER V0 ;
      RECT 2495 3335 2665 3505 ;
    LAYER V0 ;
      RECT 2495 3675 2665 3845 ;
    LAYER V0 ;
      RECT 2495 3675 2665 3845 ;
    LAYER V0 ;
      RECT 2925 3335 3095 3505 ;
    LAYER V0 ;
      RECT 2925 3675 3095 3845 ;
    LAYER V0 ;
      RECT 2925 5375 3095 5545 ;
    LAYER V0 ;
      RECT 2925 7475 3095 7645 ;
    LAYER V0 ;
      RECT 3355 3335 3525 3505 ;
    LAYER V0 ;
      RECT 3355 3675 3525 3845 ;
  END
END DP_NMOS_B_83449181_X1_Y1
