MACRO CCP_PMOS_B_53083828_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CCP_PMOS_B_53083828_X1_Y1 0 0 ;
  SIZE 5160 BY 9240 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 7420 3180 7700 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2010 1100 2290 5620 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2440 1520 2720 6040 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1550 1960 3610 2240 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 2025 1175 2275 4705 ;
    LAYER M1 ;
      RECT 2025 4955 2275 5965 ;
    LAYER M1 ;
      RECT 2025 7055 2275 8065 ;
    LAYER M1 ;
      RECT 1595 1175 1845 4705 ;
    LAYER M1 ;
      RECT 2455 1175 2705 4705 ;
    LAYER M1 ;
      RECT 2885 1175 3135 4705 ;
    LAYER M1 ;
      RECT 2885 4955 3135 5965 ;
    LAYER M1 ;
      RECT 2885 7055 3135 8065 ;
    LAYER M1 ;
      RECT 3315 1175 3565 4705 ;
    LAYER M2 ;
      RECT 1120 1120 2320 1400 ;
    LAYER M2 ;
      RECT 1980 5320 3180 5600 ;
    LAYER M2 ;
      RECT 1980 1540 3180 1820 ;
    LAYER M2 ;
      RECT 1550 5740 2750 6020 ;
    LAYER V1 ;
      RECT 2065 1175 2235 1345 ;
    LAYER V1 ;
      RECT 2065 5795 2235 5965 ;
    LAYER V1 ;
      RECT 2065 7475 2235 7645 ;
    LAYER V1 ;
      RECT 2925 1595 3095 1765 ;
    LAYER V1 ;
      RECT 2925 5375 3095 5545 ;
    LAYER V1 ;
      RECT 2925 7475 3095 7645 ;
    LAYER V1 ;
      RECT 1635 2015 1805 2185 ;
    LAYER V1 ;
      RECT 2495 2015 2665 2185 ;
    LAYER V1 ;
      RECT 3355 2015 3525 2185 ;
    LAYER V2 ;
      RECT 2075 1185 2225 1335 ;
    LAYER V2 ;
      RECT 2075 5385 2225 5535 ;
    LAYER V2 ;
      RECT 2505 1605 2655 1755 ;
    LAYER V2 ;
      RECT 2505 5805 2655 5955 ;
    LAYER V0 ;
      RECT 2065 3545 2235 3715 ;
    LAYER V0 ;
      RECT 2065 5375 2235 5545 ;
    LAYER V0 ;
      RECT 2065 7475 2235 7645 ;
    LAYER V0 ;
      RECT 1635 3545 1805 3715 ;
    LAYER V0 ;
      RECT 2495 3545 2665 3715 ;
    LAYER V0 ;
      RECT 2495 3545 2665 3715 ;
    LAYER V0 ;
      RECT 2925 3545 3095 3715 ;
    LAYER V0 ;
      RECT 2925 5375 3095 5545 ;
    LAYER V0 ;
      RECT 2925 7475 3095 7645 ;
    LAYER V0 ;
      RECT 3355 3545 3525 3715 ;
  END
END CCP_PMOS_B_53083828_X1_Y1
MACRO DP_PMOS_B_25364157_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DP_PMOS_B_25364157_X1_Y1 0 0 ;
  SIZE 5160 BY 9240 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 7420 3180 7700 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 1120 2320 1400 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 1540 3180 1820 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 5320 2320 5600 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 5740 3180 6020 ;
    END
  END GB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1550 1960 3610 2240 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 2025 1175 2275 4705 ;
    LAYER M1 ;
      RECT 2025 4955 2275 5965 ;
    LAYER M1 ;
      RECT 2025 7055 2275 8065 ;
    LAYER M1 ;
      RECT 1595 1175 1845 4705 ;
    LAYER M1 ;
      RECT 2455 1175 2705 4705 ;
    LAYER M1 ;
      RECT 2885 1175 3135 4705 ;
    LAYER M1 ;
      RECT 2885 4955 3135 5965 ;
    LAYER M1 ;
      RECT 2885 7055 3135 8065 ;
    LAYER M1 ;
      RECT 3315 1175 3565 4705 ;
    LAYER V1 ;
      RECT 2065 1175 2235 1345 ;
    LAYER V1 ;
      RECT 2065 5375 2235 5545 ;
    LAYER V1 ;
      RECT 2065 7475 2235 7645 ;
    LAYER V1 ;
      RECT 2925 1595 3095 1765 ;
    LAYER V1 ;
      RECT 2925 5795 3095 5965 ;
    LAYER V1 ;
      RECT 2925 7475 3095 7645 ;
    LAYER V1 ;
      RECT 1635 2015 1805 2185 ;
    LAYER V1 ;
      RECT 2495 2015 2665 2185 ;
    LAYER V1 ;
      RECT 3355 2015 3525 2185 ;
    LAYER V0 ;
      RECT 2065 3125 2235 3295 ;
    LAYER V0 ;
      RECT 2065 3465 2235 3635 ;
    LAYER V0 ;
      RECT 2065 3805 2235 3975 ;
    LAYER V0 ;
      RECT 2065 5375 2235 5545 ;
    LAYER V0 ;
      RECT 2065 7475 2235 7645 ;
    LAYER V0 ;
      RECT 1635 3125 1805 3295 ;
    LAYER V0 ;
      RECT 1635 3465 1805 3635 ;
    LAYER V0 ;
      RECT 1635 3805 1805 3975 ;
    LAYER V0 ;
      RECT 2495 3125 2665 3295 ;
    LAYER V0 ;
      RECT 2495 3125 2665 3295 ;
    LAYER V0 ;
      RECT 2495 3465 2665 3635 ;
    LAYER V0 ;
      RECT 2495 3465 2665 3635 ;
    LAYER V0 ;
      RECT 2495 3805 2665 3975 ;
    LAYER V0 ;
      RECT 2495 3805 2665 3975 ;
    LAYER V0 ;
      RECT 2925 3125 3095 3295 ;
    LAYER V0 ;
      RECT 2925 3465 3095 3635 ;
    LAYER V0 ;
      RECT 2925 3805 3095 3975 ;
    LAYER V0 ;
      RECT 2925 5375 3095 5545 ;
    LAYER V0 ;
      RECT 2925 7475 3095 7645 ;
    LAYER V0 ;
      RECT 3355 3125 3525 3295 ;
    LAYER V0 ;
      RECT 3355 3465 3525 3635 ;
    LAYER V0 ;
      RECT 3355 3805 3525 3975 ;
  END
END DP_PMOS_B_25364157_X1_Y1
MACRO DCAP_PMOS_57222488_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DCAP_PMOS_57222488_X1_Y1 0 0 ;
  SIZE 15480 BY 9240 ;
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6710 5320 7910 5600 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 8030 1100 8310 7720 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 7615 1175 7865 4705 ;
    LAYER M1 ;
      RECT 7615 4955 7865 5965 ;
    LAYER M1 ;
      RECT 7615 7055 7865 8065 ;
    LAYER M1 ;
      RECT 1595 1175 1845 4705 ;
    LAYER M1 ;
      RECT 13635 1175 13885 4705 ;
    LAYER M2 ;
      RECT 7140 7420 8340 7700 ;
    LAYER M2 ;
      RECT 7140 1120 8340 1400 ;
    LAYER M2 ;
      RECT 1550 1540 13930 1820 ;
    LAYER V1 ;
      RECT 7655 1175 7825 1345 ;
    LAYER V1 ;
      RECT 7655 5375 7825 5545 ;
    LAYER V1 ;
      RECT 7655 7475 7825 7645 ;
    LAYER V1 ;
      RECT 1635 1595 1805 1765 ;
    LAYER V1 ;
      RECT 13675 1595 13845 1765 ;
    LAYER V2 ;
      RECT 8095 1185 8245 1335 ;
    LAYER V2 ;
      RECT 8095 1605 8245 1755 ;
    LAYER V2 ;
      RECT 8095 7485 8245 7635 ;
    LAYER V0 ;
      RECT 7655 2705 7825 2875 ;
    LAYER V0 ;
      RECT 7655 3045 7825 3215 ;
    LAYER V0 ;
      RECT 7655 3385 7825 3555 ;
    LAYER V0 ;
      RECT 7655 3725 7825 3895 ;
    LAYER V0 ;
      RECT 7655 4065 7825 4235 ;
    LAYER V0 ;
      RECT 7655 5375 7825 5545 ;
    LAYER V0 ;
      RECT 7655 7475 7825 7645 ;
    LAYER V0 ;
      RECT 1635 2705 1805 2875 ;
    LAYER V0 ;
      RECT 1635 3045 1805 3215 ;
    LAYER V0 ;
      RECT 1635 3385 1805 3555 ;
    LAYER V0 ;
      RECT 1635 3725 1805 3895 ;
    LAYER V0 ;
      RECT 1635 4065 1805 4235 ;
    LAYER V0 ;
      RECT 13675 2705 13845 2875 ;
    LAYER V0 ;
      RECT 13675 3045 13845 3215 ;
    LAYER V0 ;
      RECT 13675 3385 13845 3555 ;
    LAYER V0 ;
      RECT 13675 3725 13845 3895 ;
    LAYER V0 ;
      RECT 13675 4065 13845 4235 ;
  END
END DCAP_PMOS_57222488_X1_Y1
MACRO CCP_NMOS_B_26073270_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CCP_NMOS_B_26073270_X1_Y1 0 0 ;
  SIZE 5160 BY 9240 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 7420 3180 7700 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2010 1100 2290 5620 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2440 1520 2720 6040 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1550 1960 3610 2240 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 2025 1175 2275 4705 ;
    LAYER M1 ;
      RECT 2025 4955 2275 5965 ;
    LAYER M1 ;
      RECT 2025 7055 2275 8065 ;
    LAYER M1 ;
      RECT 1595 1175 1845 4705 ;
    LAYER M1 ;
      RECT 2455 1175 2705 4705 ;
    LAYER M1 ;
      RECT 2885 1175 3135 4705 ;
    LAYER M1 ;
      RECT 2885 4955 3135 5965 ;
    LAYER M1 ;
      RECT 2885 7055 3135 8065 ;
    LAYER M1 ;
      RECT 3315 1175 3565 4705 ;
    LAYER M2 ;
      RECT 1120 1120 2320 1400 ;
    LAYER M2 ;
      RECT 1980 5320 3180 5600 ;
    LAYER M2 ;
      RECT 1980 1540 3180 1820 ;
    LAYER M2 ;
      RECT 1550 5740 2750 6020 ;
    LAYER V1 ;
      RECT 2065 1175 2235 1345 ;
    LAYER V1 ;
      RECT 2065 5795 2235 5965 ;
    LAYER V1 ;
      RECT 2065 7475 2235 7645 ;
    LAYER V1 ;
      RECT 2925 1595 3095 1765 ;
    LAYER V1 ;
      RECT 2925 5375 3095 5545 ;
    LAYER V1 ;
      RECT 2925 7475 3095 7645 ;
    LAYER V1 ;
      RECT 1635 2015 1805 2185 ;
    LAYER V1 ;
      RECT 2495 2015 2665 2185 ;
    LAYER V1 ;
      RECT 3355 2015 3525 2185 ;
    LAYER V2 ;
      RECT 2075 1185 2225 1335 ;
    LAYER V2 ;
      RECT 2075 5385 2225 5535 ;
    LAYER V2 ;
      RECT 2505 1605 2655 1755 ;
    LAYER V2 ;
      RECT 2505 5805 2655 5955 ;
    LAYER V0 ;
      RECT 2065 3545 2235 3715 ;
    LAYER V0 ;
      RECT 2065 5375 2235 5545 ;
    LAYER V0 ;
      RECT 2065 7475 2235 7645 ;
    LAYER V0 ;
      RECT 1635 3545 1805 3715 ;
    LAYER V0 ;
      RECT 2495 3545 2665 3715 ;
    LAYER V0 ;
      RECT 2495 3545 2665 3715 ;
    LAYER V0 ;
      RECT 2925 3545 3095 3715 ;
    LAYER V0 ;
      RECT 2925 5375 3095 5545 ;
    LAYER V0 ;
      RECT 2925 7475 3095 7645 ;
    LAYER V0 ;
      RECT 3355 3545 3525 3715 ;
  END
END CCP_NMOS_B_26073270_X1_Y1
MACRO DP_NMOS_B_83449181_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_83449181_X1_Y1 0 0 ;
  SIZE 5160 BY 9240 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 7420 3180 7700 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 1120 2320 1400 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 1540 3180 1820 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 5320 2320 5600 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 5740 3180 6020 ;
    END
  END GB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1550 1960 3610 2240 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 2025 1175 2275 4705 ;
    LAYER M1 ;
      RECT 2025 4955 2275 5965 ;
    LAYER M1 ;
      RECT 2025 7055 2275 8065 ;
    LAYER M1 ;
      RECT 1595 1175 1845 4705 ;
    LAYER M1 ;
      RECT 2455 1175 2705 4705 ;
    LAYER M1 ;
      RECT 2885 1175 3135 4705 ;
    LAYER M1 ;
      RECT 2885 4955 3135 5965 ;
    LAYER M1 ;
      RECT 2885 7055 3135 8065 ;
    LAYER M1 ;
      RECT 3315 1175 3565 4705 ;
    LAYER V1 ;
      RECT 2065 1175 2235 1345 ;
    LAYER V1 ;
      RECT 2065 5375 2235 5545 ;
    LAYER V1 ;
      RECT 2065 7475 2235 7645 ;
    LAYER V1 ;
      RECT 2925 1595 3095 1765 ;
    LAYER V1 ;
      RECT 2925 5795 3095 5965 ;
    LAYER V1 ;
      RECT 2925 7475 3095 7645 ;
    LAYER V1 ;
      RECT 1635 2015 1805 2185 ;
    LAYER V1 ;
      RECT 2495 2015 2665 2185 ;
    LAYER V1 ;
      RECT 3355 2015 3525 2185 ;
    LAYER V0 ;
      RECT 2065 3335 2235 3505 ;
    LAYER V0 ;
      RECT 2065 3675 2235 3845 ;
    LAYER V0 ;
      RECT 2065 5375 2235 5545 ;
    LAYER V0 ;
      RECT 2065 7475 2235 7645 ;
    LAYER V0 ;
      RECT 1635 3335 1805 3505 ;
    LAYER V0 ;
      RECT 1635 3675 1805 3845 ;
    LAYER V0 ;
      RECT 2495 3335 2665 3505 ;
    LAYER V0 ;
      RECT 2495 3335 2665 3505 ;
    LAYER V0 ;
      RECT 2495 3675 2665 3845 ;
    LAYER V0 ;
      RECT 2495 3675 2665 3845 ;
    LAYER V0 ;
      RECT 2925 3335 3095 3505 ;
    LAYER V0 ;
      RECT 2925 3675 3095 3845 ;
    LAYER V0 ;
      RECT 2925 5375 3095 5545 ;
    LAYER V0 ;
      RECT 2925 7475 3095 7645 ;
    LAYER V0 ;
      RECT 3355 3335 3525 3505 ;
    LAYER V0 ;
      RECT 3355 3675 3525 3845 ;
  END
END DP_NMOS_B_83449181_X1_Y1
