* power mux: DCDC_MUX
.subckt DCDC_MUX_PMOS VPWR SEL SEL_INV VIN VOUT
M1  VIN SEL_INV VOUT VPWR sky130_fd_pr__pfet_01v8 w=1050e-9 l=150e-9 nf=6 m=1
M2  VOUT SEL VIN VPWR sky130_fd_pr__pfet_01v8 w=1050e-9 l=150e-9 nf=6 m=1
.ends DCDC_MUX_PMOS

.subckt DCDC_MUX_NMOS VGND SEL SEL_INV VIN VOUT
M1  VIN SEL_INV VOUT VGND sky130_fd_pr__nfet_01v8 w=1050e-9 l=150e-9 nf=6 m=1
M2  VOUT SEL VIN VGND sky130_fd_pr__nfet_01v8 w=1050e-9 l=150e-9 nf=6 m=1
.ends DCDC_MUX_NMOS

.subckt DCDC_MUX_TGATE VGND VPWR SEL SEL_INV VIN VOUT
M1  VOUT SEL_INV VIN VPWR sky130_fd_pr__pfet_01v8 w=1050e-9 l=150e-9 nf=6 m=1
M2  VOUT SEL VIN VGND sky130_fd_pr__nfet_01v8 w=1050e-9 l=150e-9 nf=6 m=1
.ends DCDC_MUX_TGATE

.subckt inv_4 A VGND VNB VPB VPWR Y
M1 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=1050e-9 l=150e-9 nf=2 m=1
M2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1050e-9 l=150e-9 nf=4 m=1
.ends inv_4

.subckt DCDC_MUX VGND VPWR SEL_H SEL_L VIN VOUT_H VOUT_L
x0 SEL_H VGND VGND VPWR VPWR SEL_INV_H inv_4
x1 SEL_L VGND VGND VPWR VPWR SEL_INV_L inv_4
* Top MUX rail
x2 VPWR SEL_INV_H SEL_INV_H VPWR VOUT_H DCDC_MUX_PMOS
* Top MUX mid
x3 VGND VPWR SEL_INV_H SEL_H VIN VOUT_H DCDC_MUX_TGATE
* Bot MUX mid
x4 VGND VPWR SEL_L SEL_INV_L VIN VOUT_L DCDC_MUX_TGATE
* Bot MUX rail
x5 VGND SEL_INV_L SEL_INV_L VGND VOUT_L DCDC_MUX_NMOS
.ends DCDC_MUX