MACRO DCDC_CONV2TO1_1
  ORIGIN 0 0 ;
  FOREIGN DCDC_CONV2TO1_1 0 0 ;
  SIZE 72.24 BY 36.96 ;
  PIN CLK0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 7.17 19.58 7.45 26.2 ;
      LAYER M3 ;
        RECT 64.79 19.58 65.07 26.2 ;
      LAYER M3 ;
        RECT 7.17 22.495 7.45 22.865 ;
      LAYER M2 ;
        RECT 7.31 22.54 64.93 22.82 ;
      LAYER M3 ;
        RECT 64.79 22.495 65.07 22.865 ;
    END
  END CLK0
  PIN CLK0B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 28.67 10.76 28.95 17.38 ;
      LAYER M3 ;
        RECT 43.29 10.76 43.57 17.38 ;
      LAYER M3 ;
        RECT 28.67 13.675 28.95 14.045 ;
      LAYER M2 ;
        RECT 28.81 13.72 43.43 14 ;
      LAYER M3 ;
        RECT 43.29 13.675 43.57 14.045 ;
    END
  END CLK0B
  PIN CLK1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 28.67 19.58 28.95 26.2 ;
      LAYER M3 ;
        RECT 43.29 19.58 43.57 26.2 ;
      LAYER M3 ;
        RECT 28.67 22.495 28.95 22.865 ;
      LAYER M4 ;
        RECT 28.81 22.28 43.43 23.08 ;
      LAYER M3 ;
        RECT 43.29 22.495 43.57 22.865 ;
    END
  END CLK1
  PIN CLK1B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 7.17 10.76 7.45 17.38 ;
      LAYER M3 ;
        RECT 64.79 10.76 65.07 17.38 ;
      LAYER M3 ;
        RECT 7.17 13.675 7.45 14.045 ;
      LAYER M4 ;
        RECT 7.31 13.46 64.93 14.26 ;
      LAYER M3 ;
        RECT 64.79 13.675 65.07 14.045 ;
    END
  END CLK1B
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 17.46 35.14 18.66 35.42 ;
      LAYER M2 ;
        RECT 17.46 25.9 18.66 26.18 ;
      LAYER M2 ;
        RECT 17.47 35.14 17.79 35.42 ;
      LAYER M3 ;
        RECT 17.49 26.04 17.77 35.28 ;
      LAYER M2 ;
        RECT 17.47 25.9 17.79 26.18 ;
      LAYER M2 ;
        RECT 53.58 35.14 54.78 35.42 ;
      LAYER M2 ;
        RECT 53.58 25.9 54.78 26.18 ;
      LAYER M2 ;
        RECT 54.45 35.14 54.77 35.42 ;
      LAYER M3 ;
        RECT 54.47 26.04 54.75 35.28 ;
      LAYER M2 ;
        RECT 54.45 25.9 54.77 26.18 ;
      LAYER M2 ;
        RECT 18.49 35.14 53.75 35.42 ;
    END
  END VGND
  PIN VHIGH
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 17.03 7 19.09 7.28 ;
      LAYER M2 ;
        RECT 17.03 16.24 19.09 16.52 ;
      LAYER M2 ;
        RECT 17.04 7 17.36 7.28 ;
      LAYER M3 ;
        RECT 17.06 7.14 17.34 16.38 ;
      LAYER M2 ;
        RECT 17.04 16.24 17.36 16.52 ;
    END
  END VHIGH
  PIN VMID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 17.03 29.68 19.09 29.96 ;
      LAYER M2 ;
        RECT 17.03 20.44 19.09 20.72 ;
      LAYER M2 ;
        RECT 17.04 29.68 17.36 29.96 ;
      LAYER M3 ;
        RECT 17.06 20.58 17.34 29.82 ;
      LAYER M2 ;
        RECT 17.04 20.44 17.36 20.72 ;
      LAYER M2 ;
        RECT 53.15 7 55.21 7.28 ;
      LAYER M2 ;
        RECT 53.15 16.24 55.21 16.52 ;
      LAYER M2 ;
        RECT 54.88 7 55.2 7.28 ;
      LAYER M3 ;
        RECT 54.9 7.14 55.18 16.38 ;
      LAYER M2 ;
        RECT 54.88 16.24 55.2 16.52 ;
      LAYER M2 ;
        RECT 18.92 20.44 19.78 20.72 ;
      LAYER M1 ;
        RECT 19.655 16.38 19.905 20.58 ;
      LAYER M2 ;
        RECT 19.78 16.24 53.32 16.52 ;
    END
  END VMID
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 17.46 1.54 18.66 1.82 ;
      LAYER M2 ;
        RECT 17.46 10.78 18.66 11.06 ;
      LAYER M2 ;
        RECT 17.47 1.54 17.79 1.82 ;
      LAYER M3 ;
        RECT 17.49 1.68 17.77 10.92 ;
      LAYER M2 ;
        RECT 17.47 10.78 17.79 11.06 ;
      LAYER M2 ;
        RECT 53.58 1.54 54.78 1.82 ;
      LAYER M2 ;
        RECT 53.58 10.78 54.78 11.06 ;
      LAYER M2 ;
        RECT 54.45 1.54 54.77 1.82 ;
      LAYER M3 ;
        RECT 54.47 1.68 54.75 10.92 ;
      LAYER M2 ;
        RECT 54.45 10.78 54.77 11.06 ;
      LAYER M2 ;
        RECT 18.49 1.54 53.75 1.82 ;
    END
  END VPWR
  PIN Y0_TOP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 18.32 17.08 19.52 17.36 ;
      LAYER M2 ;
        RECT 18.32 19.6 19.52 19.88 ;
      LAYER M2 ;
        RECT 18.76 17.08 19.08 17.36 ;
      LAYER M3 ;
        RECT 18.78 17.22 19.06 19.74 ;
      LAYER M2 ;
        RECT 18.76 19.6 19.08 19.88 ;
    END
  END Y0_TOP
  PIN Y1_TOP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 17.46 16.66 18.66 16.94 ;
      LAYER M2 ;
        RECT 17.46 20.02 18.66 20.3 ;
      LAYER M2 ;
        RECT 17.9 16.66 18.22 16.94 ;
      LAYER M3 ;
        RECT 17.92 16.8 18.2 20.16 ;
      LAYER M2 ;
        RECT 17.9 20.02 18.22 20.3 ;
    END
  END Y1_TOP
  PIN VLOW
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 53.15 29.68 55.21 29.96 ;
      LAYER M2 ;
        RECT 53.15 20.44 55.21 20.72 ;
      LAYER M2 ;
        RECT 54.88 29.68 55.2 29.96 ;
      LAYER M3 ;
        RECT 54.9 20.58 55.18 29.82 ;
      LAYER M2 ;
        RECT 54.88 20.44 55.2 20.72 ;
    END
  END VLOW
  PIN Y0_BOT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 52.72 17.08 53.92 17.36 ;
      LAYER M2 ;
        RECT 52.72 19.6 53.92 19.88 ;
      LAYER M2 ;
        RECT 53.16 17.08 53.48 17.36 ;
      LAYER M3 ;
        RECT 53.18 17.22 53.46 19.74 ;
      LAYER M2 ;
        RECT 53.16 19.6 53.48 19.88 ;
    END
  END Y0_BOT
  PIN Y1_BOT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 53.58 16.66 54.78 16.94 ;
      LAYER M2 ;
        RECT 53.58 20.02 54.78 20.3 ;
      LAYER M2 ;
        RECT 54.02 16.66 54.34 16.94 ;
      LAYER M3 ;
        RECT 54.04 16.8 54.32 20.16 ;
      LAYER M2 ;
        RECT 54.02 20.02 54.34 20.3 ;
    END
  END Y1_BOT
  OBS 
  LAYER M3 ;
        RECT 18.35 3.62 18.63 8.14 ;
  LAYER M2 ;
        RECT 18.32 12.88 19.52 13.16 ;
  LAYER M2 ;
        RECT 27.35 12.88 28.55 13.16 ;
  LAYER M3 ;
        RECT 18.35 7.98 18.63 13.02 ;
  LAYER M2 ;
        RECT 18.33 12.88 18.65 13.16 ;
  LAYER M2 ;
        RECT 19.35 12.88 27.52 13.16 ;
  LAYER M2 ;
        RECT 18.33 12.88 18.65 13.16 ;
  LAYER M3 ;
        RECT 18.35 12.86 18.63 13.18 ;
  LAYER M2 ;
        RECT 18.33 12.88 18.65 13.16 ;
  LAYER M3 ;
        RECT 18.35 12.86 18.63 13.18 ;
  LAYER M2 ;
        RECT 18.33 12.88 18.65 13.16 ;
  LAYER M3 ;
        RECT 18.35 12.86 18.63 13.18 ;
  LAYER M2 ;
        RECT 18.33 12.88 18.65 13.16 ;
  LAYER M3 ;
        RECT 18.35 12.86 18.63 13.18 ;
  LAYER M3 ;
        RECT 17.92 3.2 18.2 7.72 ;
  LAYER M2 ;
        RECT 17.46 12.46 18.66 12.74 ;
  LAYER M2 ;
        RECT 7.57 12.88 8.77 13.16 ;
  LAYER M3 ;
        RECT 17.92 7.56 18.2 12.6 ;
  LAYER M2 ;
        RECT 17.9 12.46 18.22 12.74 ;
  LAYER M2 ;
        RECT 17.47 12.46 17.79 12.74 ;
  LAYER M3 ;
        RECT 17.49 12.6 17.77 13.02 ;
  LAYER M2 ;
        RECT 8.6 12.88 17.63 13.16 ;
  LAYER M2 ;
        RECT 17.9 12.46 18.22 12.74 ;
  LAYER M3 ;
        RECT 17.92 12.44 18.2 12.76 ;
  LAYER M2 ;
        RECT 17.9 12.46 18.22 12.74 ;
  LAYER M3 ;
        RECT 17.92 12.44 18.2 12.76 ;
  LAYER M2 ;
        RECT 17.47 12.46 17.79 12.74 ;
  LAYER M3 ;
        RECT 17.49 12.44 17.77 12.76 ;
  LAYER M2 ;
        RECT 17.47 12.88 17.79 13.16 ;
  LAYER M3 ;
        RECT 17.49 12.86 17.77 13.18 ;
  LAYER M2 ;
        RECT 17.9 12.46 18.22 12.74 ;
  LAYER M3 ;
        RECT 17.92 12.44 18.2 12.76 ;
  LAYER M2 ;
        RECT 17.47 12.46 17.79 12.74 ;
  LAYER M3 ;
        RECT 17.49 12.44 17.77 12.76 ;
  LAYER M2 ;
        RECT 17.47 12.88 17.79 13.16 ;
  LAYER M3 ;
        RECT 17.49 12.86 17.77 13.18 ;
  LAYER M2 ;
        RECT 17.9 12.46 18.22 12.74 ;
  LAYER M3 ;
        RECT 17.92 12.44 18.2 12.76 ;
  LAYER M1 ;
        RECT 18.365 4.535 18.615 8.065 ;
  LAYER M1 ;
        RECT 18.365 3.275 18.615 4.285 ;
  LAYER M1 ;
        RECT 18.365 1.175 18.615 2.185 ;
  LAYER M1 ;
        RECT 18.795 4.535 19.045 8.065 ;
  LAYER M1 ;
        RECT 17.935 4.535 18.185 8.065 ;
  LAYER M1 ;
        RECT 17.505 4.535 17.755 8.065 ;
  LAYER M1 ;
        RECT 17.505 3.275 17.755 4.285 ;
  LAYER M1 ;
        RECT 17.505 1.175 17.755 2.185 ;
  LAYER M1 ;
        RECT 17.075 4.535 17.325 8.065 ;
  LAYER M2 ;
        RECT 18.32 7.84 19.52 8.12 ;
  LAYER M2 ;
        RECT 17.46 3.64 18.66 3.92 ;
  LAYER M2 ;
        RECT 17.46 7.42 18.66 7.7 ;
  LAYER M2 ;
        RECT 17.89 3.22 19.09 3.5 ;
  LAYER M2 ;
        RECT 17.46 1.54 18.66 1.82 ;
  LAYER M3 ;
        RECT 18.35 3.62 18.63 8.14 ;
  LAYER M3 ;
        RECT 17.92 3.2 18.2 7.72 ;
  LAYER M2 ;
        RECT 17.03 7 19.09 7.28 ;
  LAYER M1 ;
        RECT 18.365 13.775 18.615 17.305 ;
  LAYER M1 ;
        RECT 18.365 12.515 18.615 13.525 ;
  LAYER M1 ;
        RECT 18.365 10.415 18.615 11.425 ;
  LAYER M1 ;
        RECT 18.795 13.775 19.045 17.305 ;
  LAYER M1 ;
        RECT 17.935 13.775 18.185 17.305 ;
  LAYER M1 ;
        RECT 17.505 13.775 17.755 17.305 ;
  LAYER M1 ;
        RECT 17.505 12.515 17.755 13.525 ;
  LAYER M1 ;
        RECT 17.505 10.415 17.755 11.425 ;
  LAYER M1 ;
        RECT 17.075 13.775 17.325 17.305 ;
  LAYER M2 ;
        RECT 17.46 10.78 18.66 11.06 ;
  LAYER M2 ;
        RECT 18.32 17.08 19.52 17.36 ;
  LAYER M2 ;
        RECT 17.46 16.66 18.66 16.94 ;
  LAYER M2 ;
        RECT 18.32 12.88 19.52 13.16 ;
  LAYER M2 ;
        RECT 17.46 12.46 18.66 12.74 ;
  LAYER M2 ;
        RECT 17.03 16.24 19.09 16.52 ;
  LAYER M1 ;
        RECT 28.255 13.775 28.505 17.305 ;
  LAYER M1 ;
        RECT 28.255 12.515 28.505 13.525 ;
  LAYER M1 ;
        RECT 28.255 10.415 28.505 11.425 ;
  LAYER M1 ;
        RECT 22.235 13.775 22.485 17.305 ;
  LAYER M1 ;
        RECT 34.275 13.775 34.525 17.305 ;
  LAYER M2 ;
        RECT 27.78 10.78 28.98 11.06 ;
  LAYER M2 ;
        RECT 27.78 17.08 28.98 17.36 ;
  LAYER M2 ;
        RECT 22.19 16.66 34.57 16.94 ;
  LAYER M2 ;
        RECT 27.35 12.88 28.55 13.16 ;
  LAYER M3 ;
        RECT 28.67 10.76 28.95 17.38 ;
  LAYER M1 ;
        RECT 7.615 13.775 7.865 17.305 ;
  LAYER M1 ;
        RECT 7.615 12.515 7.865 13.525 ;
  LAYER M1 ;
        RECT 7.615 10.415 7.865 11.425 ;
  LAYER M1 ;
        RECT 13.635 13.775 13.885 17.305 ;
  LAYER M1 ;
        RECT 1.595 13.775 1.845 17.305 ;
  LAYER M2 ;
        RECT 7.14 10.78 8.34 11.06 ;
  LAYER M2 ;
        RECT 7.14 17.08 8.34 17.36 ;
  LAYER M2 ;
        RECT 1.55 16.66 13.93 16.94 ;
  LAYER M2 ;
        RECT 7.57 12.88 8.77 13.16 ;
  LAYER M3 ;
        RECT 7.17 10.76 7.45 17.38 ;
  LAYER M3 ;
        RECT 18.35 28.82 18.63 33.34 ;
  LAYER M2 ;
        RECT 18.32 23.8 19.52 24.08 ;
  LAYER M2 ;
        RECT 27.35 23.8 28.55 24.08 ;
  LAYER M3 ;
        RECT 18.35 23.94 18.63 28.98 ;
  LAYER M2 ;
        RECT 18.33 23.8 18.65 24.08 ;
  LAYER M2 ;
        RECT 19.35 23.8 27.52 24.08 ;
  LAYER M2 ;
        RECT 18.33 23.8 18.65 24.08 ;
  LAYER M3 ;
        RECT 18.35 23.78 18.63 24.1 ;
  LAYER M2 ;
        RECT 18.33 23.8 18.65 24.08 ;
  LAYER M3 ;
        RECT 18.35 23.78 18.63 24.1 ;
  LAYER M2 ;
        RECT 18.33 23.8 18.65 24.08 ;
  LAYER M3 ;
        RECT 18.35 23.78 18.63 24.1 ;
  LAYER M2 ;
        RECT 18.33 23.8 18.65 24.08 ;
  LAYER M3 ;
        RECT 18.35 23.78 18.63 24.1 ;
  LAYER M3 ;
        RECT 17.92 29.24 18.2 33.76 ;
  LAYER M2 ;
        RECT 17.46 24.22 18.66 24.5 ;
  LAYER M2 ;
        RECT 7.57 23.8 8.77 24.08 ;
  LAYER M3 ;
        RECT 17.92 24.36 18.2 29.4 ;
  LAYER M2 ;
        RECT 17.9 24.22 18.22 24.5 ;
  LAYER M2 ;
        RECT 17.47 24.22 17.79 24.5 ;
  LAYER M3 ;
        RECT 17.49 23.94 17.77 24.36 ;
  LAYER M2 ;
        RECT 8.6 23.8 17.63 24.08 ;
  LAYER M2 ;
        RECT 17.9 24.22 18.22 24.5 ;
  LAYER M3 ;
        RECT 17.92 24.2 18.2 24.52 ;
  LAYER M2 ;
        RECT 17.9 24.22 18.22 24.5 ;
  LAYER M3 ;
        RECT 17.92 24.2 18.2 24.52 ;
  LAYER M2 ;
        RECT 17.47 24.22 17.79 24.5 ;
  LAYER M3 ;
        RECT 17.49 24.2 17.77 24.52 ;
  LAYER M2 ;
        RECT 17.47 23.8 17.79 24.08 ;
  LAYER M3 ;
        RECT 17.49 23.78 17.77 24.1 ;
  LAYER M2 ;
        RECT 17.9 24.22 18.22 24.5 ;
  LAYER M3 ;
        RECT 17.92 24.2 18.2 24.52 ;
  LAYER M2 ;
        RECT 17.47 24.22 17.79 24.5 ;
  LAYER M3 ;
        RECT 17.49 24.2 17.77 24.52 ;
  LAYER M2 ;
        RECT 17.47 23.8 17.79 24.08 ;
  LAYER M3 ;
        RECT 17.49 23.78 17.77 24.1 ;
  LAYER M2 ;
        RECT 17.9 24.22 18.22 24.5 ;
  LAYER M3 ;
        RECT 17.92 24.2 18.2 24.52 ;
  LAYER M1 ;
        RECT 18.365 28.895 18.615 32.425 ;
  LAYER M1 ;
        RECT 18.365 32.675 18.615 33.685 ;
  LAYER M1 ;
        RECT 18.365 34.775 18.615 35.785 ;
  LAYER M1 ;
        RECT 18.795 28.895 19.045 32.425 ;
  LAYER M1 ;
        RECT 17.935 28.895 18.185 32.425 ;
  LAYER M1 ;
        RECT 17.505 28.895 17.755 32.425 ;
  LAYER M1 ;
        RECT 17.505 32.675 17.755 33.685 ;
  LAYER M1 ;
        RECT 17.505 34.775 17.755 35.785 ;
  LAYER M1 ;
        RECT 17.075 28.895 17.325 32.425 ;
  LAYER M2 ;
        RECT 18.32 28.84 19.52 29.12 ;
  LAYER M2 ;
        RECT 17.46 33.04 18.66 33.32 ;
  LAYER M2 ;
        RECT 17.46 29.26 18.66 29.54 ;
  LAYER M2 ;
        RECT 17.89 33.46 19.09 33.74 ;
  LAYER M2 ;
        RECT 17.46 35.14 18.66 35.42 ;
  LAYER M3 ;
        RECT 18.35 28.82 18.63 33.34 ;
  LAYER M3 ;
        RECT 17.92 29.24 18.2 33.76 ;
  LAYER M2 ;
        RECT 17.03 29.68 19.09 29.96 ;
  LAYER M1 ;
        RECT 18.365 19.655 18.615 23.185 ;
  LAYER M1 ;
        RECT 18.365 23.435 18.615 24.445 ;
  LAYER M1 ;
        RECT 18.365 25.535 18.615 26.545 ;
  LAYER M1 ;
        RECT 18.795 19.655 19.045 23.185 ;
  LAYER M1 ;
        RECT 17.935 19.655 18.185 23.185 ;
  LAYER M1 ;
        RECT 17.505 19.655 17.755 23.185 ;
  LAYER M1 ;
        RECT 17.505 23.435 17.755 24.445 ;
  LAYER M1 ;
        RECT 17.505 25.535 17.755 26.545 ;
  LAYER M1 ;
        RECT 17.075 19.655 17.325 23.185 ;
  LAYER M2 ;
        RECT 17.46 25.9 18.66 26.18 ;
  LAYER M2 ;
        RECT 18.32 19.6 19.52 19.88 ;
  LAYER M2 ;
        RECT 17.46 20.02 18.66 20.3 ;
  LAYER M2 ;
        RECT 18.32 23.8 19.52 24.08 ;
  LAYER M2 ;
        RECT 17.46 24.22 18.66 24.5 ;
  LAYER M2 ;
        RECT 17.03 20.44 19.09 20.72 ;
  LAYER M1 ;
        RECT 28.255 19.655 28.505 23.185 ;
  LAYER M1 ;
        RECT 28.255 23.435 28.505 24.445 ;
  LAYER M1 ;
        RECT 28.255 25.535 28.505 26.545 ;
  LAYER M1 ;
        RECT 22.235 19.655 22.485 23.185 ;
  LAYER M1 ;
        RECT 34.275 19.655 34.525 23.185 ;
  LAYER M2 ;
        RECT 27.78 25.9 28.98 26.18 ;
  LAYER M2 ;
        RECT 27.78 19.6 28.98 19.88 ;
  LAYER M2 ;
        RECT 22.19 20.02 34.57 20.3 ;
  LAYER M2 ;
        RECT 27.35 23.8 28.55 24.08 ;
  LAYER M3 ;
        RECT 28.67 19.58 28.95 26.2 ;
  LAYER M1 ;
        RECT 7.615 19.655 7.865 23.185 ;
  LAYER M1 ;
        RECT 7.615 23.435 7.865 24.445 ;
  LAYER M1 ;
        RECT 7.615 25.535 7.865 26.545 ;
  LAYER M1 ;
        RECT 13.635 19.655 13.885 23.185 ;
  LAYER M1 ;
        RECT 1.595 19.655 1.845 23.185 ;
  LAYER M2 ;
        RECT 7.14 25.9 8.34 26.18 ;
  LAYER M2 ;
        RECT 7.14 19.6 8.34 19.88 ;
  LAYER M2 ;
        RECT 1.55 20.02 13.93 20.3 ;
  LAYER M2 ;
        RECT 7.57 23.8 8.77 24.08 ;
  LAYER M3 ;
        RECT 7.17 19.58 7.45 26.2 ;
  LAYER M3 ;
        RECT 53.61 3.62 53.89 8.14 ;
  LAYER M2 ;
        RECT 52.72 12.88 53.92 13.16 ;
  LAYER M2 ;
        RECT 43.69 12.88 44.89 13.16 ;
  LAYER M3 ;
        RECT 53.61 7.98 53.89 13.02 ;
  LAYER M2 ;
        RECT 53.59 12.88 53.91 13.16 ;
  LAYER M2 ;
        RECT 44.72 12.88 52.89 13.16 ;
  LAYER M2 ;
        RECT 53.59 12.88 53.91 13.16 ;
  LAYER M3 ;
        RECT 53.61 12.86 53.89 13.18 ;
  LAYER M2 ;
        RECT 53.59 12.88 53.91 13.16 ;
  LAYER M3 ;
        RECT 53.61 12.86 53.89 13.18 ;
  LAYER M2 ;
        RECT 53.59 12.88 53.91 13.16 ;
  LAYER M3 ;
        RECT 53.61 12.86 53.89 13.18 ;
  LAYER M2 ;
        RECT 53.59 12.88 53.91 13.16 ;
  LAYER M3 ;
        RECT 53.61 12.86 53.89 13.18 ;
  LAYER M3 ;
        RECT 54.04 3.2 54.32 7.72 ;
  LAYER M2 ;
        RECT 53.58 12.46 54.78 12.74 ;
  LAYER M2 ;
        RECT 63.47 12.88 64.67 13.16 ;
  LAYER M3 ;
        RECT 54.04 7.56 54.32 12.6 ;
  LAYER M2 ;
        RECT 54.02 12.46 54.34 12.74 ;
  LAYER M2 ;
        RECT 54.45 12.46 54.77 12.74 ;
  LAYER M3 ;
        RECT 54.47 12.6 54.75 13.02 ;
  LAYER M2 ;
        RECT 54.61 12.88 63.64 13.16 ;
  LAYER M2 ;
        RECT 54.02 12.46 54.34 12.74 ;
  LAYER M3 ;
        RECT 54.04 12.44 54.32 12.76 ;
  LAYER M2 ;
        RECT 54.02 12.46 54.34 12.74 ;
  LAYER M3 ;
        RECT 54.04 12.44 54.32 12.76 ;
  LAYER M2 ;
        RECT 54.45 12.46 54.77 12.74 ;
  LAYER M3 ;
        RECT 54.47 12.44 54.75 12.76 ;
  LAYER M2 ;
        RECT 54.45 12.88 54.77 13.16 ;
  LAYER M3 ;
        RECT 54.47 12.86 54.75 13.18 ;
  LAYER M2 ;
        RECT 54.02 12.46 54.34 12.74 ;
  LAYER M3 ;
        RECT 54.04 12.44 54.32 12.76 ;
  LAYER M2 ;
        RECT 54.45 12.46 54.77 12.74 ;
  LAYER M3 ;
        RECT 54.47 12.44 54.75 12.76 ;
  LAYER M2 ;
        RECT 54.45 12.88 54.77 13.16 ;
  LAYER M3 ;
        RECT 54.47 12.86 54.75 13.18 ;
  LAYER M2 ;
        RECT 54.02 12.46 54.34 12.74 ;
  LAYER M3 ;
        RECT 54.04 12.44 54.32 12.76 ;
  LAYER M1 ;
        RECT 53.625 4.535 53.875 8.065 ;
  LAYER M1 ;
        RECT 53.625 3.275 53.875 4.285 ;
  LAYER M1 ;
        RECT 53.625 1.175 53.875 2.185 ;
  LAYER M1 ;
        RECT 53.195 4.535 53.445 8.065 ;
  LAYER M1 ;
        RECT 54.055 4.535 54.305 8.065 ;
  LAYER M1 ;
        RECT 54.485 4.535 54.735 8.065 ;
  LAYER M1 ;
        RECT 54.485 3.275 54.735 4.285 ;
  LAYER M1 ;
        RECT 54.485 1.175 54.735 2.185 ;
  LAYER M1 ;
        RECT 54.915 4.535 55.165 8.065 ;
  LAYER M2 ;
        RECT 52.72 7.84 53.92 8.12 ;
  LAYER M2 ;
        RECT 53.58 3.64 54.78 3.92 ;
  LAYER M2 ;
        RECT 53.58 7.42 54.78 7.7 ;
  LAYER M2 ;
        RECT 53.15 3.22 54.35 3.5 ;
  LAYER M2 ;
        RECT 53.58 1.54 54.78 1.82 ;
  LAYER M3 ;
        RECT 53.61 3.62 53.89 8.14 ;
  LAYER M3 ;
        RECT 54.04 3.2 54.32 7.72 ;
  LAYER M2 ;
        RECT 53.15 7 55.21 7.28 ;
  LAYER M1 ;
        RECT 53.625 13.775 53.875 17.305 ;
  LAYER M1 ;
        RECT 53.625 12.515 53.875 13.525 ;
  LAYER M1 ;
        RECT 53.625 10.415 53.875 11.425 ;
  LAYER M1 ;
        RECT 53.195 13.775 53.445 17.305 ;
  LAYER M1 ;
        RECT 54.055 13.775 54.305 17.305 ;
  LAYER M1 ;
        RECT 54.485 13.775 54.735 17.305 ;
  LAYER M1 ;
        RECT 54.485 12.515 54.735 13.525 ;
  LAYER M1 ;
        RECT 54.485 10.415 54.735 11.425 ;
  LAYER M1 ;
        RECT 54.915 13.775 55.165 17.305 ;
  LAYER M2 ;
        RECT 53.58 10.78 54.78 11.06 ;
  LAYER M2 ;
        RECT 52.72 17.08 53.92 17.36 ;
  LAYER M2 ;
        RECT 53.58 16.66 54.78 16.94 ;
  LAYER M2 ;
        RECT 52.72 12.88 53.92 13.16 ;
  LAYER M2 ;
        RECT 53.58 12.46 54.78 12.74 ;
  LAYER M2 ;
        RECT 53.15 16.24 55.21 16.52 ;
  LAYER M1 ;
        RECT 43.735 13.775 43.985 17.305 ;
  LAYER M1 ;
        RECT 43.735 12.515 43.985 13.525 ;
  LAYER M1 ;
        RECT 43.735 10.415 43.985 11.425 ;
  LAYER M1 ;
        RECT 49.755 13.775 50.005 17.305 ;
  LAYER M1 ;
        RECT 37.715 13.775 37.965 17.305 ;
  LAYER M2 ;
        RECT 43.26 10.78 44.46 11.06 ;
  LAYER M2 ;
        RECT 43.26 17.08 44.46 17.36 ;
  LAYER M2 ;
        RECT 37.67 16.66 50.05 16.94 ;
  LAYER M2 ;
        RECT 43.69 12.88 44.89 13.16 ;
  LAYER M3 ;
        RECT 43.29 10.76 43.57 17.38 ;
  LAYER M1 ;
        RECT 64.375 13.775 64.625 17.305 ;
  LAYER M1 ;
        RECT 64.375 12.515 64.625 13.525 ;
  LAYER M1 ;
        RECT 64.375 10.415 64.625 11.425 ;
  LAYER M1 ;
        RECT 58.355 13.775 58.605 17.305 ;
  LAYER M1 ;
        RECT 70.395 13.775 70.645 17.305 ;
  LAYER M2 ;
        RECT 63.9 10.78 65.1 11.06 ;
  LAYER M2 ;
        RECT 63.9 17.08 65.1 17.36 ;
  LAYER M2 ;
        RECT 58.31 16.66 70.69 16.94 ;
  LAYER M2 ;
        RECT 63.47 12.88 64.67 13.16 ;
  LAYER M3 ;
        RECT 64.79 10.76 65.07 17.38 ;
  LAYER M3 ;
        RECT 53.61 28.82 53.89 33.34 ;
  LAYER M2 ;
        RECT 52.72 23.8 53.92 24.08 ;
  LAYER M2 ;
        RECT 43.69 23.8 44.89 24.08 ;
  LAYER M3 ;
        RECT 53.61 23.94 53.89 28.98 ;
  LAYER M2 ;
        RECT 53.59 23.8 53.91 24.08 ;
  LAYER M2 ;
        RECT 44.72 23.8 52.89 24.08 ;
  LAYER M2 ;
        RECT 53.59 23.8 53.91 24.08 ;
  LAYER M3 ;
        RECT 53.61 23.78 53.89 24.1 ;
  LAYER M2 ;
        RECT 53.59 23.8 53.91 24.08 ;
  LAYER M3 ;
        RECT 53.61 23.78 53.89 24.1 ;
  LAYER M2 ;
        RECT 53.59 23.8 53.91 24.08 ;
  LAYER M3 ;
        RECT 53.61 23.78 53.89 24.1 ;
  LAYER M2 ;
        RECT 53.59 23.8 53.91 24.08 ;
  LAYER M3 ;
        RECT 53.61 23.78 53.89 24.1 ;
  LAYER M3 ;
        RECT 54.04 29.24 54.32 33.76 ;
  LAYER M2 ;
        RECT 53.58 24.22 54.78 24.5 ;
  LAYER M2 ;
        RECT 63.47 23.8 64.67 24.08 ;
  LAYER M3 ;
        RECT 54.04 24.36 54.32 29.4 ;
  LAYER M2 ;
        RECT 54.02 24.22 54.34 24.5 ;
  LAYER M2 ;
        RECT 54.45 24.22 54.77 24.5 ;
  LAYER M3 ;
        RECT 54.47 23.94 54.75 24.36 ;
  LAYER M2 ;
        RECT 54.61 23.8 63.64 24.08 ;
  LAYER M2 ;
        RECT 54.02 24.22 54.34 24.5 ;
  LAYER M3 ;
        RECT 54.04 24.2 54.32 24.52 ;
  LAYER M2 ;
        RECT 54.02 24.22 54.34 24.5 ;
  LAYER M3 ;
        RECT 54.04 24.2 54.32 24.52 ;
  LAYER M2 ;
        RECT 54.45 24.22 54.77 24.5 ;
  LAYER M3 ;
        RECT 54.47 24.2 54.75 24.52 ;
  LAYER M2 ;
        RECT 54.45 23.8 54.77 24.08 ;
  LAYER M3 ;
        RECT 54.47 23.78 54.75 24.1 ;
  LAYER M2 ;
        RECT 54.02 24.22 54.34 24.5 ;
  LAYER M3 ;
        RECT 54.04 24.2 54.32 24.52 ;
  LAYER M2 ;
        RECT 54.45 24.22 54.77 24.5 ;
  LAYER M3 ;
        RECT 54.47 24.2 54.75 24.52 ;
  LAYER M2 ;
        RECT 54.45 23.8 54.77 24.08 ;
  LAYER M3 ;
        RECT 54.47 23.78 54.75 24.1 ;
  LAYER M2 ;
        RECT 54.02 24.22 54.34 24.5 ;
  LAYER M3 ;
        RECT 54.04 24.2 54.32 24.52 ;
  LAYER M1 ;
        RECT 53.625 28.895 53.875 32.425 ;
  LAYER M1 ;
        RECT 53.625 32.675 53.875 33.685 ;
  LAYER M1 ;
        RECT 53.625 34.775 53.875 35.785 ;
  LAYER M1 ;
        RECT 53.195 28.895 53.445 32.425 ;
  LAYER M1 ;
        RECT 54.055 28.895 54.305 32.425 ;
  LAYER M1 ;
        RECT 54.485 28.895 54.735 32.425 ;
  LAYER M1 ;
        RECT 54.485 32.675 54.735 33.685 ;
  LAYER M1 ;
        RECT 54.485 34.775 54.735 35.785 ;
  LAYER M1 ;
        RECT 54.915 28.895 55.165 32.425 ;
  LAYER M2 ;
        RECT 52.72 28.84 53.92 29.12 ;
  LAYER M2 ;
        RECT 53.58 33.04 54.78 33.32 ;
  LAYER M2 ;
        RECT 53.58 29.26 54.78 29.54 ;
  LAYER M2 ;
        RECT 53.15 33.46 54.35 33.74 ;
  LAYER M2 ;
        RECT 53.58 35.14 54.78 35.42 ;
  LAYER M3 ;
        RECT 53.61 28.82 53.89 33.34 ;
  LAYER M3 ;
        RECT 54.04 29.24 54.32 33.76 ;
  LAYER M2 ;
        RECT 53.15 29.68 55.21 29.96 ;
  LAYER M1 ;
        RECT 53.625 19.655 53.875 23.185 ;
  LAYER M1 ;
        RECT 53.625 23.435 53.875 24.445 ;
  LAYER M1 ;
        RECT 53.625 25.535 53.875 26.545 ;
  LAYER M1 ;
        RECT 53.195 19.655 53.445 23.185 ;
  LAYER M1 ;
        RECT 54.055 19.655 54.305 23.185 ;
  LAYER M1 ;
        RECT 54.485 19.655 54.735 23.185 ;
  LAYER M1 ;
        RECT 54.485 23.435 54.735 24.445 ;
  LAYER M1 ;
        RECT 54.485 25.535 54.735 26.545 ;
  LAYER M1 ;
        RECT 54.915 19.655 55.165 23.185 ;
  LAYER M2 ;
        RECT 53.58 25.9 54.78 26.18 ;
  LAYER M2 ;
        RECT 52.72 19.6 53.92 19.88 ;
  LAYER M2 ;
        RECT 53.58 20.02 54.78 20.3 ;
  LAYER M2 ;
        RECT 52.72 23.8 53.92 24.08 ;
  LAYER M2 ;
        RECT 53.58 24.22 54.78 24.5 ;
  LAYER M2 ;
        RECT 53.15 20.44 55.21 20.72 ;
  LAYER M1 ;
        RECT 43.735 19.655 43.985 23.185 ;
  LAYER M1 ;
        RECT 43.735 23.435 43.985 24.445 ;
  LAYER M1 ;
        RECT 43.735 25.535 43.985 26.545 ;
  LAYER M1 ;
        RECT 49.755 19.655 50.005 23.185 ;
  LAYER M1 ;
        RECT 37.715 19.655 37.965 23.185 ;
  LAYER M2 ;
        RECT 43.26 25.9 44.46 26.18 ;
  LAYER M2 ;
        RECT 43.26 19.6 44.46 19.88 ;
  LAYER M2 ;
        RECT 37.67 20.02 50.05 20.3 ;
  LAYER M2 ;
        RECT 43.69 23.8 44.89 24.08 ;
  LAYER M3 ;
        RECT 43.29 19.58 43.57 26.2 ;
  LAYER M1 ;
        RECT 64.375 19.655 64.625 23.185 ;
  LAYER M1 ;
        RECT 64.375 23.435 64.625 24.445 ;
  LAYER M1 ;
        RECT 64.375 25.535 64.625 26.545 ;
  LAYER M1 ;
        RECT 58.355 19.655 58.605 23.185 ;
  LAYER M1 ;
        RECT 70.395 19.655 70.645 23.185 ;
  LAYER M2 ;
        RECT 63.9 25.9 65.1 26.18 ;
  LAYER M2 ;
        RECT 63.9 19.6 65.1 19.88 ;
  LAYER M2 ;
        RECT 58.31 20.02 70.69 20.3 ;
  LAYER M2 ;
        RECT 63.47 23.8 64.67 24.08 ;
  LAYER M3 ;
        RECT 64.79 19.58 65.07 26.2 ;
  END 
END DCDC_CONV2TO1_1
