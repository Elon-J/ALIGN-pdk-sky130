MACRO CAP_2T_55207366
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CAP_2T_55207366 0 0 ;
  SIZE 1000001980 BY 1000005300 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 265 860 1000001285 1660 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 265 1000003640 1000001285 1000004440 ;
    END
  END PLUS
  OBS
    LAYER M4 ;
      RECT 860 2370 1000001160 1000002670 ;
    LAYER M4 ;
      RECT 1000000710 1000001320 1000001160 1000003840 ;
    LAYER M5 ;
      RECT 1085 830 1535 3350 ;
    LAYER V4 ;
      RECT 1210 1160 1410 1360 ;
  END
END CAP_2T_55207366
