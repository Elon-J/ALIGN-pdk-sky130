MACRO DCDC_XSW_PMOS
  ORIGIN 0 0 ;
  FOREIGN DCDC_XSW_PMOS 0 0 ;
  SIZE 36.12 BY 18.48 ;
  PIN VPB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 17.46 16.66 18.66 16.94 ;
      LAYER M2 ;
        RECT 17.46 7.42 18.66 7.7 ;
      LAYER M2 ;
        RECT 17.47 16.66 17.79 16.94 ;
      LAYER M3 ;
        RECT 17.49 7.56 17.77 16.8 ;
      LAYER M2 ;
        RECT 17.47 7.42 17.79 7.7 ;
    END
  END VPB
  PIN VIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 17.03 11.2 19.09 11.48 ;
      LAYER M2 ;
        RECT 17.03 1.96 19.09 2.24 ;
      LAYER M2 ;
        RECT 17.04 11.2 17.36 11.48 ;
      LAYER M3 ;
        RECT 17.06 2.1 17.34 11.34 ;
      LAYER M2 ;
        RECT 17.04 1.96 17.36 2.24 ;
    END
  END VIN
  PIN VOUT0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 18.32 1.12 19.52 1.4 ;
    END
  END VOUT0
  PIN VOUT1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 17.46 1.54 18.66 1.82 ;
    END
  END VOUT1
  PIN CLKB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 28.67 1.1 28.95 7.72 ;
    END
  END CLKB
  PIN CLK
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 7.17 1.1 7.45 7.72 ;
    END
  END CLK
  OBS 
  LAYER M3 ;
        RECT 18.35 10.34 18.63 14.86 ;
  LAYER M2 ;
        RECT 18.32 5.32 19.52 5.6 ;
  LAYER M2 ;
        RECT 27.35 5.32 28.55 5.6 ;
  LAYER M3 ;
        RECT 18.35 5.46 18.63 10.5 ;
  LAYER M2 ;
        RECT 18.33 5.32 18.65 5.6 ;
  LAYER M2 ;
        RECT 19.35 5.32 27.52 5.6 ;
  LAYER M2 ;
        RECT 18.33 5.32 18.65 5.6 ;
  LAYER M3 ;
        RECT 18.35 5.3 18.63 5.62 ;
  LAYER M2 ;
        RECT 18.33 5.32 18.65 5.6 ;
  LAYER M3 ;
        RECT 18.35 5.3 18.63 5.62 ;
  LAYER M2 ;
        RECT 18.33 5.32 18.65 5.6 ;
  LAYER M3 ;
        RECT 18.35 5.3 18.63 5.62 ;
  LAYER M2 ;
        RECT 18.33 5.32 18.65 5.6 ;
  LAYER M3 ;
        RECT 18.35 5.3 18.63 5.62 ;
  LAYER M3 ;
        RECT 17.92 10.76 18.2 15.28 ;
  LAYER M2 ;
        RECT 17.46 5.74 18.66 6.02 ;
  LAYER M2 ;
        RECT 7.57 5.32 8.77 5.6 ;
  LAYER M3 ;
        RECT 17.92 5.88 18.2 10.92 ;
  LAYER M2 ;
        RECT 17.9 5.74 18.22 6.02 ;
  LAYER M2 ;
        RECT 17.47 5.74 17.79 6.02 ;
  LAYER M3 ;
        RECT 17.49 5.46 17.77 5.88 ;
  LAYER M2 ;
        RECT 8.6 5.32 17.63 5.6 ;
  LAYER M2 ;
        RECT 17.9 5.74 18.22 6.02 ;
  LAYER M3 ;
        RECT 17.92 5.72 18.2 6.04 ;
  LAYER M2 ;
        RECT 17.9 5.74 18.22 6.02 ;
  LAYER M3 ;
        RECT 17.92 5.72 18.2 6.04 ;
  LAYER M2 ;
        RECT 17.47 5.74 17.79 6.02 ;
  LAYER M3 ;
        RECT 17.49 5.72 17.77 6.04 ;
  LAYER M2 ;
        RECT 17.47 5.32 17.79 5.6 ;
  LAYER M3 ;
        RECT 17.49 5.3 17.77 5.62 ;
  LAYER M2 ;
        RECT 17.9 5.74 18.22 6.02 ;
  LAYER M3 ;
        RECT 17.92 5.72 18.2 6.04 ;
  LAYER M2 ;
        RECT 17.47 5.74 17.79 6.02 ;
  LAYER M3 ;
        RECT 17.49 5.72 17.77 6.04 ;
  LAYER M2 ;
        RECT 17.47 5.32 17.79 5.6 ;
  LAYER M3 ;
        RECT 17.49 5.3 17.77 5.62 ;
  LAYER M2 ;
        RECT 17.9 5.74 18.22 6.02 ;
  LAYER M3 ;
        RECT 17.92 5.72 18.2 6.04 ;
  LAYER M1 ;
        RECT 18.365 10.415 18.615 13.945 ;
  LAYER M1 ;
        RECT 18.365 14.195 18.615 15.205 ;
  LAYER M1 ;
        RECT 18.365 16.295 18.615 17.305 ;
  LAYER M1 ;
        RECT 18.795 10.415 19.045 13.945 ;
  LAYER M1 ;
        RECT 17.935 10.415 18.185 13.945 ;
  LAYER M1 ;
        RECT 17.505 10.415 17.755 13.945 ;
  LAYER M1 ;
        RECT 17.505 14.195 17.755 15.205 ;
  LAYER M1 ;
        RECT 17.505 16.295 17.755 17.305 ;
  LAYER M1 ;
        RECT 17.075 10.415 17.325 13.945 ;
  LAYER M2 ;
        RECT 17.46 14.56 18.66 14.84 ;
  LAYER M2 ;
        RECT 18.32 10.36 19.52 10.64 ;
  LAYER M2 ;
        RECT 17.89 14.98 19.09 15.26 ;
  LAYER M2 ;
        RECT 17.46 10.78 18.66 11.06 ;
  LAYER M2 ;
        RECT 17.46 16.66 18.66 16.94 ;
  LAYER M3 ;
        RECT 18.35 10.34 18.63 14.86 ;
  LAYER M3 ;
        RECT 17.92 10.76 18.2 15.28 ;
  LAYER M2 ;
        RECT 17.03 11.2 19.09 11.48 ;
  LAYER M1 ;
        RECT 18.365 1.175 18.615 4.705 ;
  LAYER M1 ;
        RECT 18.365 4.955 18.615 5.965 ;
  LAYER M1 ;
        RECT 18.365 7.055 18.615 8.065 ;
  LAYER M1 ;
        RECT 18.795 1.175 19.045 4.705 ;
  LAYER M1 ;
        RECT 17.935 1.175 18.185 4.705 ;
  LAYER M1 ;
        RECT 17.505 1.175 17.755 4.705 ;
  LAYER M1 ;
        RECT 17.505 4.955 17.755 5.965 ;
  LAYER M1 ;
        RECT 17.505 7.055 17.755 8.065 ;
  LAYER M1 ;
        RECT 17.075 1.175 17.325 4.705 ;
  LAYER M2 ;
        RECT 17.46 7.42 18.66 7.7 ;
  LAYER M2 ;
        RECT 18.32 1.12 19.52 1.4 ;
  LAYER M2 ;
        RECT 17.46 1.54 18.66 1.82 ;
  LAYER M2 ;
        RECT 18.32 5.32 19.52 5.6 ;
  LAYER M2 ;
        RECT 17.46 5.74 18.66 6.02 ;
  LAYER M2 ;
        RECT 17.03 1.96 19.09 2.24 ;
  LAYER M1 ;
        RECT 28.255 1.175 28.505 4.705 ;
  LAYER M1 ;
        RECT 28.255 4.955 28.505 5.965 ;
  LAYER M1 ;
        RECT 28.255 7.055 28.505 8.065 ;
  LAYER M1 ;
        RECT 22.235 1.175 22.485 4.705 ;
  LAYER M1 ;
        RECT 34.275 1.175 34.525 4.705 ;
  LAYER M2 ;
        RECT 22.19 1.12 34.57 1.4 ;
  LAYER M2 ;
        RECT 27.78 7.42 28.98 7.7 ;
  LAYER M2 ;
        RECT 27.78 1.54 28.98 1.82 ;
  LAYER M2 ;
        RECT 27.35 5.32 28.55 5.6 ;
  LAYER M3 ;
        RECT 28.67 1.1 28.95 7.72 ;
  LAYER M1 ;
        RECT 7.615 1.175 7.865 4.705 ;
  LAYER M1 ;
        RECT 7.615 4.955 7.865 5.965 ;
  LAYER M1 ;
        RECT 7.615 7.055 7.865 8.065 ;
  LAYER M1 ;
        RECT 13.635 1.175 13.885 4.705 ;
  LAYER M1 ;
        RECT 1.595 1.175 1.845 4.705 ;
  LAYER M2 ;
        RECT 1.55 1.12 13.93 1.4 ;
  LAYER M2 ;
        RECT 7.14 7.42 8.34 7.7 ;
  LAYER M2 ;
        RECT 7.14 1.54 8.34 1.82 ;
  LAYER M2 ;
        RECT 7.57 5.32 8.77 5.6 ;
  LAYER M3 ;
        RECT 7.17 1.1 7.45 7.72 ;
  END 
END DCDC_XSW_PMOS
