MACRO DCDC_XSW_NMOS
  ORIGIN 0 0 ;
  FOREIGN DCDC_XSW_NMOS 0 0 ;
  SIZE 36.12 BY 18.48 ;
  PIN VNB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 17.46 1.54 18.66 1.82 ;
      LAYER M2 ;
        RECT 17.46 10.78 18.66 11.06 ;
      LAYER M2 ;
        RECT 17.47 1.54 17.79 1.82 ;
      LAYER M3 ;
        RECT 17.49 1.68 17.77 10.92 ;
      LAYER M2 ;
        RECT 17.47 10.78 17.79 11.06 ;
    END
  END VNB
  PIN VIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 17.03 7 19.09 7.28 ;
      LAYER M2 ;
        RECT 17.03 16.24 19.09 16.52 ;
      LAYER M2 ;
        RECT 17.04 7 17.36 7.28 ;
      LAYER M3 ;
        RECT 17.06 7.14 17.34 16.38 ;
      LAYER M2 ;
        RECT 17.04 16.24 17.36 16.52 ;
    END
  END VIN
  PIN VOUT0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 18.32 17.08 19.52 17.36 ;
    END
  END VOUT0
  PIN VOUT1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 17.46 16.66 18.66 16.94 ;
    END
  END VOUT1
  PIN CLKB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 28.67 10.76 28.95 17.38 ;
    END
  END CLKB
  PIN CLK
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 7.17 10.76 7.45 17.38 ;
    END
  END CLK
  OBS 
  LAYER M3 ;
        RECT 18.35 3.62 18.63 8.14 ;
  LAYER M2 ;
        RECT 18.32 12.88 19.52 13.16 ;
  LAYER M2 ;
        RECT 27.35 12.88 28.55 13.16 ;
  LAYER M3 ;
        RECT 18.35 7.98 18.63 13.02 ;
  LAYER M2 ;
        RECT 18.33 12.88 18.65 13.16 ;
  LAYER M2 ;
        RECT 19.35 12.88 27.52 13.16 ;
  LAYER M2 ;
        RECT 18.33 12.88 18.65 13.16 ;
  LAYER M3 ;
        RECT 18.35 12.86 18.63 13.18 ;
  LAYER M2 ;
        RECT 18.33 12.88 18.65 13.16 ;
  LAYER M3 ;
        RECT 18.35 12.86 18.63 13.18 ;
  LAYER M2 ;
        RECT 18.33 12.88 18.65 13.16 ;
  LAYER M3 ;
        RECT 18.35 12.86 18.63 13.18 ;
  LAYER M2 ;
        RECT 18.33 12.88 18.65 13.16 ;
  LAYER M3 ;
        RECT 18.35 12.86 18.63 13.18 ;
  LAYER M3 ;
        RECT 17.92 3.2 18.2 7.72 ;
  LAYER M2 ;
        RECT 17.46 12.46 18.66 12.74 ;
  LAYER M2 ;
        RECT 7.57 12.88 8.77 13.16 ;
  LAYER M3 ;
        RECT 17.92 7.56 18.2 12.6 ;
  LAYER M2 ;
        RECT 17.9 12.46 18.22 12.74 ;
  LAYER M2 ;
        RECT 17.47 12.46 17.79 12.74 ;
  LAYER M3 ;
        RECT 17.49 12.6 17.77 13.02 ;
  LAYER M2 ;
        RECT 8.6 12.88 17.63 13.16 ;
  LAYER M2 ;
        RECT 17.9 12.46 18.22 12.74 ;
  LAYER M3 ;
        RECT 17.92 12.44 18.2 12.76 ;
  LAYER M2 ;
        RECT 17.9 12.46 18.22 12.74 ;
  LAYER M3 ;
        RECT 17.92 12.44 18.2 12.76 ;
  LAYER M2 ;
        RECT 17.47 12.46 17.79 12.74 ;
  LAYER M3 ;
        RECT 17.49 12.44 17.77 12.76 ;
  LAYER M2 ;
        RECT 17.47 12.88 17.79 13.16 ;
  LAYER M3 ;
        RECT 17.49 12.86 17.77 13.18 ;
  LAYER M2 ;
        RECT 17.9 12.46 18.22 12.74 ;
  LAYER M3 ;
        RECT 17.92 12.44 18.2 12.76 ;
  LAYER M2 ;
        RECT 17.47 12.46 17.79 12.74 ;
  LAYER M3 ;
        RECT 17.49 12.44 17.77 12.76 ;
  LAYER M2 ;
        RECT 17.47 12.88 17.79 13.16 ;
  LAYER M3 ;
        RECT 17.49 12.86 17.77 13.18 ;
  LAYER M2 ;
        RECT 17.9 12.46 18.22 12.74 ;
  LAYER M3 ;
        RECT 17.92 12.44 18.2 12.76 ;
  LAYER M1 ;
        RECT 18.365 4.535 18.615 8.065 ;
  LAYER M1 ;
        RECT 18.365 3.275 18.615 4.285 ;
  LAYER M1 ;
        RECT 18.365 1.175 18.615 2.185 ;
  LAYER M1 ;
        RECT 18.795 4.535 19.045 8.065 ;
  LAYER M1 ;
        RECT 17.935 4.535 18.185 8.065 ;
  LAYER M1 ;
        RECT 17.505 4.535 17.755 8.065 ;
  LAYER M1 ;
        RECT 17.505 3.275 17.755 4.285 ;
  LAYER M1 ;
        RECT 17.505 1.175 17.755 2.185 ;
  LAYER M1 ;
        RECT 17.075 4.535 17.325 8.065 ;
  LAYER M2 ;
        RECT 18.32 7.84 19.52 8.12 ;
  LAYER M2 ;
        RECT 17.46 3.64 18.66 3.92 ;
  LAYER M2 ;
        RECT 17.46 7.42 18.66 7.7 ;
  LAYER M2 ;
        RECT 17.89 3.22 19.09 3.5 ;
  LAYER M2 ;
        RECT 17.46 1.54 18.66 1.82 ;
  LAYER M3 ;
        RECT 18.35 3.62 18.63 8.14 ;
  LAYER M3 ;
        RECT 17.92 3.2 18.2 7.72 ;
  LAYER M2 ;
        RECT 17.03 7 19.09 7.28 ;
  LAYER M1 ;
        RECT 18.365 13.775 18.615 17.305 ;
  LAYER M1 ;
        RECT 18.365 12.515 18.615 13.525 ;
  LAYER M1 ;
        RECT 18.365 10.415 18.615 11.425 ;
  LAYER M1 ;
        RECT 18.795 13.775 19.045 17.305 ;
  LAYER M1 ;
        RECT 17.935 13.775 18.185 17.305 ;
  LAYER M1 ;
        RECT 17.505 13.775 17.755 17.305 ;
  LAYER M1 ;
        RECT 17.505 12.515 17.755 13.525 ;
  LAYER M1 ;
        RECT 17.505 10.415 17.755 11.425 ;
  LAYER M1 ;
        RECT 17.075 13.775 17.325 17.305 ;
  LAYER M2 ;
        RECT 17.46 10.78 18.66 11.06 ;
  LAYER M2 ;
        RECT 18.32 17.08 19.52 17.36 ;
  LAYER M2 ;
        RECT 17.46 16.66 18.66 16.94 ;
  LAYER M2 ;
        RECT 18.32 12.88 19.52 13.16 ;
  LAYER M2 ;
        RECT 17.46 12.46 18.66 12.74 ;
  LAYER M2 ;
        RECT 17.03 16.24 19.09 16.52 ;
  LAYER M1 ;
        RECT 28.255 13.775 28.505 17.305 ;
  LAYER M1 ;
        RECT 28.255 12.515 28.505 13.525 ;
  LAYER M1 ;
        RECT 28.255 10.415 28.505 11.425 ;
  LAYER M1 ;
        RECT 22.235 13.775 22.485 17.305 ;
  LAYER M1 ;
        RECT 34.275 13.775 34.525 17.305 ;
  LAYER M2 ;
        RECT 27.78 10.78 28.98 11.06 ;
  LAYER M2 ;
        RECT 27.78 17.08 28.98 17.36 ;
  LAYER M2 ;
        RECT 22.19 16.66 34.57 16.94 ;
  LAYER M2 ;
        RECT 27.35 12.88 28.55 13.16 ;
  LAYER M3 ;
        RECT 28.67 10.76 28.95 17.38 ;
  LAYER M1 ;
        RECT 7.615 13.775 7.865 17.305 ;
  LAYER M1 ;
        RECT 7.615 12.515 7.865 13.525 ;
  LAYER M1 ;
        RECT 7.615 10.415 7.865 11.425 ;
  LAYER M1 ;
        RECT 13.635 13.775 13.885 17.305 ;
  LAYER M1 ;
        RECT 1.595 13.775 1.845 17.305 ;
  LAYER M2 ;
        RECT 7.14 10.78 8.34 11.06 ;
  LAYER M2 ;
        RECT 7.14 17.08 8.34 17.36 ;
  LAYER M2 ;
        RECT 1.55 16.66 13.93 16.94 ;
  LAYER M2 ;
        RECT 7.57 12.88 8.77 13.16 ;
  LAYER M3 ;
        RECT 7.17 10.76 7.45 17.38 ;
  END 
END DCDC_XSW_NMOS
