* power mux: DCDC_MUX
.subckt DCDC_MUX_PMOS VPWR SEL SEL_INV VIN VOUT
m1  VIN SEL_INV VOUT VPWR sky130_fd_pr__pfet_01v8 w=2100e-9 l=150e-9 nf=2 m=3
m2  VOUT SEL     VIN VPWR sky130_fd_pr__pfet_01v8 w=2100e-9 l=150e-9 nf=2 m=3
.ends DCDC_MUX_PMOS

.subckt DCDC_MUX_NMOS VGND SEL SEL_INV VIN VOUT
m1  VIN SEL_INV VOUT VGND sky130_fd_pr__nfet_01v8 w=2100e-9 l=150e-9 nf=2 m=3
m2  VOUT SEL     VIN VGND sky130_fd_pr__nfet_01v8 w=2100e-9 l=150e-9 nf=2 m=3
.ends DCDC_MUX_NMOS

.subckt DCDC_MUX_TGATE VGND VPWR SEL SEL_INV VIN VOUT
m1  VOUT SEL_INV VIN VPWR sky130_fd_pr__pfet_01v8 w=2100e-9 l=150e-9 nf=2 m=3
m2  VOUT SEL     VIN VGND sky130_fd_pr__nfet_01v8 w=2100e-9 l=150e-9 nf=2 m=3
.ends DCDC_MUX_TGATE

.subckt DCDC_MUX VGND VPWR SEL_H SEL_INV_H SEL_L SEL_INV_L VIN VOUT_H VOUT_L
* Top MUX rail
x0 VPWR SEL_INV_H SEL_INV_H VPWR VOUT_H DCDC_MUX_PMOS
* Top MUX mid
x1 VGND VPWR SEL_INV_H SEL_H VIN VOUT_H DCDC_MUX_TGATE
* Bot MUX mid
x2 VGND VPWR SEL_L SEL_INV_L VIN VOUT_L DCDC_MUX_TGATE
* Bot MUX rail
x3 VGND SEL_INV_L SEL_INV_L VGND VOUT_L DCDC_MUX_NMOS
.ends DCDC_MUX