.subckt CAP_TEST VPWR VGND
C1 VPWR VGND sky130_fd_pr__cap_mim_m3_1 w=15 l=1
.ends CAP_TEST