MACRO CCP_PMOS_B_53083828_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CCP_PMOS_B_53083828_X1_Y1 0 0 ;
  SIZE 3440 BY 7560 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 6580 2320 6860 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1150 260 1430 4780 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 680 1860 5200 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 690 1120 2750 1400 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 7225 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M2 ;
      RECT 260 280 1460 560 ;
    LAYER M2 ;
      RECT 1120 4480 2320 4760 ;
    LAYER M2 ;
      RECT 1120 700 2320 980 ;
    LAYER M2 ;
      RECT 690 4900 1890 5180 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4955 1375 5125 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 2065 755 2235 925 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 1635 1175 1805 1345 ;
    LAYER V1 ;
      RECT 2495 1175 2665 1345 ;
    LAYER V2 ;
      RECT 1215 345 1365 495 ;
    LAYER V2 ;
      RECT 1215 4545 1365 4695 ;
    LAYER V2 ;
      RECT 1645 765 1795 915 ;
    LAYER V2 ;
      RECT 1645 4965 1795 5115 ;
    LAYER V0 ;
      RECT 1205 2705 1375 2875 ;
    LAYER V0 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V0 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V0 ;
      RECT 775 2705 945 2875 ;
    LAYER V0 ;
      RECT 1635 2705 1805 2875 ;
    LAYER V0 ;
      RECT 1635 2705 1805 2875 ;
    LAYER V0 ;
      RECT 2065 2705 2235 2875 ;
    LAYER V0 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V0 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V0 ;
      RECT 2495 2705 2665 2875 ;
  END
END CCP_PMOS_B_53083828_X1_Y1
