MACRO PMOS_4T_48942251_X1_Y2
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN PMOS_4T_48942251_X1_Y2 0 0 ;
  SIZE 4300 BY 15120 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 13300 2320 13580 ;
    END
  END B
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 1100 1860 7300 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2010 5300 2290 11500 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2440 1520 2720 7720 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 2025 1175 2275 4705 ;
    LAYER M1 ;
      RECT 2025 4955 2275 5965 ;
    LAYER M1 ;
      RECT 2025 7055 2275 10585 ;
    LAYER M1 ;
      RECT 2025 10835 2275 11845 ;
    LAYER M1 ;
      RECT 2025 12935 2275 13945 ;
    LAYER M1 ;
      RECT 1595 1175 1845 4705 ;
    LAYER M1 ;
      RECT 1595 7055 1845 10585 ;
    LAYER M1 ;
      RECT 2455 1175 2705 4705 ;
    LAYER M1 ;
      RECT 2455 7055 2705 10585 ;
    LAYER M2 ;
      RECT 1120 1120 2320 1400 ;
    LAYER M2 ;
      RECT 1120 5320 2320 5600 ;
    LAYER M2 ;
      RECT 1550 1540 2750 1820 ;
    LAYER M2 ;
      RECT 1120 7000 2320 7280 ;
    LAYER M2 ;
      RECT 1120 11200 2320 11480 ;
    LAYER M2 ;
      RECT 1550 7420 2750 7700 ;
    LAYER V1 ;
      RECT 2065 1175 2235 1345 ;
    LAYER V1 ;
      RECT 2065 5375 2235 5545 ;
    LAYER V1 ;
      RECT 2065 7055 2235 7225 ;
    LAYER V1 ;
      RECT 2065 11255 2235 11425 ;
    LAYER V1 ;
      RECT 2065 13355 2235 13525 ;
    LAYER V1 ;
      RECT 1635 1595 1805 1765 ;
    LAYER V1 ;
      RECT 1635 7475 1805 7645 ;
    LAYER V1 ;
      RECT 2495 1595 2665 1765 ;
    LAYER V1 ;
      RECT 2495 7475 2665 7645 ;
    LAYER V2 ;
      RECT 1645 1185 1795 1335 ;
    LAYER V2 ;
      RECT 1645 7065 1795 7215 ;
    LAYER V2 ;
      RECT 2075 5385 2225 5535 ;
    LAYER V2 ;
      RECT 2075 11265 2225 11415 ;
    LAYER V2 ;
      RECT 2505 1605 2655 1755 ;
    LAYER V2 ;
      RECT 2505 7485 2655 7635 ;
    LAYER V0 ;
      RECT 2065 3545 2235 3715 ;
    LAYER V0 ;
      RECT 2065 5375 2235 5545 ;
    LAYER V0 ;
      RECT 2065 9425 2235 9595 ;
    LAYER V0 ;
      RECT 2065 11255 2235 11425 ;
    LAYER V0 ;
      RECT 2065 13355 2235 13525 ;
    LAYER V0 ;
      RECT 2065 13355 2235 13525 ;
    LAYER V0 ;
      RECT 1635 3545 1805 3715 ;
    LAYER V0 ;
      RECT 1635 9425 1805 9595 ;
    LAYER V0 ;
      RECT 2495 3545 2665 3715 ;
    LAYER V0 ;
      RECT 2495 9425 2665 9595 ;
  END
END PMOS_4T_48942251_X1_Y2
