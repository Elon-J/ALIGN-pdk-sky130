MACRO DCDC_HUNIT_CONV2TO1
  ORIGIN 0 0 ;
  FOREIGN DCDC_HUNIT_CONV2TO1 0 0 ;
  SIZE 30.96 BY 30.24 ;
  PIN CLK1B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 6.31 8.24 6.59 14.86 ;
    END
  END CLK1B
  PIN CLK0B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 24.37 8.24 24.65 14.86 ;
    END
  END CLK0B
  PIN VHIGH
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.45 6.16 16.51 6.44 ;
      LAYER M2 ;
        RECT 14.45 13.72 16.51 14 ;
      LAYER M2 ;
        RECT 16.18 6.16 16.5 6.44 ;
      LAYER M3 ;
        RECT 16.2 6.3 16.48 13.86 ;
      LAYER M2 ;
        RECT 16.18 13.72 16.5 14 ;
    END
  END VHIGH
  PIN Y0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.74 14.56 16.94 14.84 ;
      LAYER M2 ;
        RECT 15.74 15.4 16.94 15.68 ;
      LAYER M2 ;
        RECT 16.18 14.56 16.5 14.84 ;
      LAYER M3 ;
        RECT 16.2 14.7 16.48 15.54 ;
      LAYER M2 ;
        RECT 16.18 15.4 16.5 15.68 ;
    END
  END Y0
  PIN Y1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.88 14.14 16.08 14.42 ;
      LAYER M2 ;
        RECT 14.88 15.82 16.08 16.1 ;
      LAYER M2 ;
        RECT 15.32 14.14 15.64 14.42 ;
      LAYER M3 ;
        RECT 15.34 14.28 15.62 15.96 ;
      LAYER M2 ;
        RECT 15.32 15.82 15.64 16.1 ;
    END
  END Y1
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.88 0.7 16.08 0.98 ;
      LAYER M2 ;
        RECT 14.88 8.26 16.08 8.54 ;
      LAYER M2 ;
        RECT 14.89 0.7 15.21 0.98 ;
      LAYER M3 ;
        RECT 14.91 0.84 15.19 8.4 ;
      LAYER M2 ;
        RECT 14.89 8.26 15.21 8.54 ;
    END
  END VPWR
  PIN CLK0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 6.31 15.38 6.59 22 ;
    END
  END CLK0
  PIN CLK1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 24.37 15.38 24.65 22 ;
    END
  END CLK1
  PIN VLOW
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.45 23.8 16.51 24.08 ;
      LAYER M2 ;
        RECT 14.45 16.24 16.51 16.52 ;
      LAYER M2 ;
        RECT 16.18 23.8 16.5 24.08 ;
      LAYER M3 ;
        RECT 16.2 16.38 16.48 23.94 ;
      LAYER M2 ;
        RECT 16.18 16.24 16.5 16.52 ;
    END
  END VLOW
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.88 29.26 16.08 29.54 ;
      LAYER M2 ;
        RECT 14.88 21.7 16.08 21.98 ;
      LAYER M2 ;
        RECT 14.89 29.26 15.21 29.54 ;
      LAYER M3 ;
        RECT 14.91 21.84 15.19 29.4 ;
      LAYER M2 ;
        RECT 14.89 21.7 15.21 21.98 ;
    END
  END VGND
  OBS 
  LAYER M3 ;
        RECT 15.77 2.78 16.05 7.3 ;
  LAYER M2 ;
        RECT 15.74 10.36 16.94 10.64 ;
  LAYER M2 ;
        RECT 23.05 10.36 24.25 10.64 ;
  LAYER M3 ;
        RECT 15.77 7.14 16.05 10.5 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M2 ;
        RECT 16.77 10.36 23.22 10.64 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M3 ;
        RECT 15.34 2.36 15.62 6.88 ;
  LAYER M2 ;
        RECT 14.88 9.94 16.08 10.22 ;
  LAYER M2 ;
        RECT 6.71 10.36 7.91 10.64 ;
  LAYER M3 ;
        RECT 15.34 6.72 15.62 10.08 ;
  LAYER M2 ;
        RECT 15.32 9.94 15.64 10.22 ;
  LAYER M2 ;
        RECT 14.89 9.94 15.21 10.22 ;
  LAYER M3 ;
        RECT 14.91 10.08 15.19 10.5 ;
  LAYER M2 ;
        RECT 7.74 10.36 15.05 10.64 ;
  LAYER M2 ;
        RECT 15.32 9.94 15.64 10.22 ;
  LAYER M3 ;
        RECT 15.34 9.92 15.62 10.24 ;
  LAYER M2 ;
        RECT 15.32 9.94 15.64 10.22 ;
  LAYER M3 ;
        RECT 15.34 9.92 15.62 10.24 ;
  LAYER M2 ;
        RECT 15.32 9.94 15.64 10.22 ;
  LAYER M3 ;
        RECT 15.34 9.92 15.62 10.24 ;
  LAYER M2 ;
        RECT 14.89 9.94 15.21 10.22 ;
  LAYER M3 ;
        RECT 14.91 9.92 15.19 10.24 ;
  LAYER M2 ;
        RECT 14.89 10.36 15.21 10.64 ;
  LAYER M3 ;
        RECT 14.91 10.34 15.19 10.66 ;
  LAYER M2 ;
        RECT 15.32 9.94 15.64 10.22 ;
  LAYER M3 ;
        RECT 15.34 9.92 15.62 10.24 ;
  LAYER M2 ;
        RECT 14.89 9.94 15.21 10.22 ;
  LAYER M3 ;
        RECT 14.91 9.92 15.19 10.24 ;
  LAYER M2 ;
        RECT 14.89 10.36 15.21 10.64 ;
  LAYER M3 ;
        RECT 14.91 10.34 15.19 10.66 ;
  LAYER M1 ;
        RECT 15.785 3.695 16.035 7.225 ;
  LAYER M1 ;
        RECT 15.785 2.435 16.035 3.445 ;
  LAYER M1 ;
        RECT 15.785 0.335 16.035 1.345 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M1 ;
        RECT 14.925 2.435 15.175 3.445 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 1.345 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M2 ;
        RECT 15.74 7 16.94 7.28 ;
  LAYER M2 ;
        RECT 14.88 2.8 16.08 3.08 ;
  LAYER M2 ;
        RECT 14.88 6.58 16.08 6.86 ;
  LAYER M2 ;
        RECT 15.31 2.38 16.51 2.66 ;
  LAYER M2 ;
        RECT 14.88 0.7 16.08 0.98 ;
  LAYER M3 ;
        RECT 15.77 2.78 16.05 7.3 ;
  LAYER M3 ;
        RECT 15.34 2.36 15.62 6.88 ;
  LAYER M2 ;
        RECT 14.45 6.16 16.51 6.44 ;
  LAYER M1 ;
        RECT 15.785 11.255 16.035 14.785 ;
  LAYER M1 ;
        RECT 15.785 9.995 16.035 11.005 ;
  LAYER M1 ;
        RECT 15.785 7.895 16.035 8.905 ;
  LAYER M1 ;
        RECT 16.215 11.255 16.465 14.785 ;
  LAYER M1 ;
        RECT 15.355 11.255 15.605 14.785 ;
  LAYER M1 ;
        RECT 14.925 11.255 15.175 14.785 ;
  LAYER M1 ;
        RECT 14.925 9.995 15.175 11.005 ;
  LAYER M1 ;
        RECT 14.925 7.895 15.175 8.905 ;
  LAYER M1 ;
        RECT 14.495 11.255 14.745 14.785 ;
  LAYER M2 ;
        RECT 14.88 8.26 16.08 8.54 ;
  LAYER M2 ;
        RECT 15.74 14.56 16.94 14.84 ;
  LAYER M2 ;
        RECT 14.88 14.14 16.08 14.42 ;
  LAYER M2 ;
        RECT 15.74 10.36 16.94 10.64 ;
  LAYER M2 ;
        RECT 14.88 9.94 16.08 10.22 ;
  LAYER M2 ;
        RECT 14.45 13.72 16.51 14 ;
  LAYER M1 ;
        RECT 23.955 11.255 24.205 14.785 ;
  LAYER M1 ;
        RECT 23.955 9.995 24.205 11.005 ;
  LAYER M1 ;
        RECT 23.955 7.895 24.205 8.905 ;
  LAYER M1 ;
        RECT 17.935 11.255 18.185 14.785 ;
  LAYER M1 ;
        RECT 29.975 11.255 30.225 14.785 ;
  LAYER M2 ;
        RECT 17.89 14.56 30.27 14.84 ;
  LAYER M2 ;
        RECT 23.48 8.26 24.68 8.54 ;
  LAYER M2 ;
        RECT 23.48 14.14 24.68 14.42 ;
  LAYER M2 ;
        RECT 23.05 10.36 24.25 10.64 ;
  LAYER M3 ;
        RECT 24.37 8.24 24.65 14.86 ;
  LAYER M1 ;
        RECT 6.755 11.255 7.005 14.785 ;
  LAYER M1 ;
        RECT 6.755 9.995 7.005 11.005 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 8.905 ;
  LAYER M1 ;
        RECT 12.775 11.255 13.025 14.785 ;
  LAYER M1 ;
        RECT 0.735 11.255 0.985 14.785 ;
  LAYER M2 ;
        RECT 0.69 14.56 13.07 14.84 ;
  LAYER M2 ;
        RECT 6.28 8.26 7.48 8.54 ;
  LAYER M2 ;
        RECT 6.28 14.14 7.48 14.42 ;
  LAYER M2 ;
        RECT 6.71 10.36 7.91 10.64 ;
  LAYER M3 ;
        RECT 6.31 8.24 6.59 14.86 ;
  LAYER M3 ;
        RECT 15.77 22.94 16.05 27.46 ;
  LAYER M2 ;
        RECT 15.74 19.6 16.94 19.88 ;
  LAYER M2 ;
        RECT 23.05 19.6 24.25 19.88 ;
  LAYER M3 ;
        RECT 15.77 19.74 16.05 23.1 ;
  LAYER M2 ;
        RECT 15.75 19.6 16.07 19.88 ;
  LAYER M2 ;
        RECT 16.77 19.6 23.22 19.88 ;
  LAYER M2 ;
        RECT 15.75 19.6 16.07 19.88 ;
  LAYER M3 ;
        RECT 15.77 19.58 16.05 19.9 ;
  LAYER M2 ;
        RECT 15.75 19.6 16.07 19.88 ;
  LAYER M3 ;
        RECT 15.77 19.58 16.05 19.9 ;
  LAYER M2 ;
        RECT 15.75 19.6 16.07 19.88 ;
  LAYER M3 ;
        RECT 15.77 19.58 16.05 19.9 ;
  LAYER M2 ;
        RECT 15.75 19.6 16.07 19.88 ;
  LAYER M3 ;
        RECT 15.77 19.58 16.05 19.9 ;
  LAYER M3 ;
        RECT 15.34 23.36 15.62 27.88 ;
  LAYER M2 ;
        RECT 14.88 20.02 16.08 20.3 ;
  LAYER M2 ;
        RECT 6.71 19.6 7.91 19.88 ;
  LAYER M3 ;
        RECT 15.34 20.16 15.62 23.52 ;
  LAYER M2 ;
        RECT 15.32 20.02 15.64 20.3 ;
  LAYER M2 ;
        RECT 14.89 20.02 15.21 20.3 ;
  LAYER M3 ;
        RECT 14.91 19.74 15.19 20.16 ;
  LAYER M2 ;
        RECT 7.74 19.6 15.05 19.88 ;
  LAYER M2 ;
        RECT 15.32 20.02 15.64 20.3 ;
  LAYER M3 ;
        RECT 15.34 20 15.62 20.32 ;
  LAYER M2 ;
        RECT 15.32 20.02 15.64 20.3 ;
  LAYER M3 ;
        RECT 15.34 20 15.62 20.32 ;
  LAYER M2 ;
        RECT 15.32 20.02 15.64 20.3 ;
  LAYER M3 ;
        RECT 15.34 20 15.62 20.32 ;
  LAYER M2 ;
        RECT 14.89 19.6 15.21 19.88 ;
  LAYER M3 ;
        RECT 14.91 19.58 15.19 19.9 ;
  LAYER M2 ;
        RECT 14.89 20.02 15.21 20.3 ;
  LAYER M3 ;
        RECT 14.91 20 15.19 20.32 ;
  LAYER M2 ;
        RECT 15.32 20.02 15.64 20.3 ;
  LAYER M3 ;
        RECT 15.34 20 15.62 20.32 ;
  LAYER M2 ;
        RECT 14.89 19.6 15.21 19.88 ;
  LAYER M3 ;
        RECT 14.91 19.58 15.19 19.9 ;
  LAYER M2 ;
        RECT 14.89 20.02 15.21 20.3 ;
  LAYER M3 ;
        RECT 14.91 20 15.19 20.32 ;
  LAYER M1 ;
        RECT 15.785 23.015 16.035 26.545 ;
  LAYER M1 ;
        RECT 15.785 26.795 16.035 27.805 ;
  LAYER M1 ;
        RECT 15.785 28.895 16.035 29.905 ;
  LAYER M1 ;
        RECT 16.215 23.015 16.465 26.545 ;
  LAYER M1 ;
        RECT 15.355 23.015 15.605 26.545 ;
  LAYER M1 ;
        RECT 14.925 23.015 15.175 26.545 ;
  LAYER M1 ;
        RECT 14.925 26.795 15.175 27.805 ;
  LAYER M1 ;
        RECT 14.925 28.895 15.175 29.905 ;
  LAYER M1 ;
        RECT 14.495 23.015 14.745 26.545 ;
  LAYER M2 ;
        RECT 15.74 22.96 16.94 23.24 ;
  LAYER M2 ;
        RECT 14.88 27.16 16.08 27.44 ;
  LAYER M2 ;
        RECT 14.88 23.38 16.08 23.66 ;
  LAYER M2 ;
        RECT 15.31 27.58 16.51 27.86 ;
  LAYER M2 ;
        RECT 14.88 29.26 16.08 29.54 ;
  LAYER M3 ;
        RECT 15.77 22.94 16.05 27.46 ;
  LAYER M3 ;
        RECT 15.34 23.36 15.62 27.88 ;
  LAYER M2 ;
        RECT 14.45 23.8 16.51 24.08 ;
  LAYER M1 ;
        RECT 15.785 15.455 16.035 18.985 ;
  LAYER M1 ;
        RECT 15.785 19.235 16.035 20.245 ;
  LAYER M1 ;
        RECT 15.785 21.335 16.035 22.345 ;
  LAYER M1 ;
        RECT 16.215 15.455 16.465 18.985 ;
  LAYER M1 ;
        RECT 15.355 15.455 15.605 18.985 ;
  LAYER M1 ;
        RECT 14.925 15.455 15.175 18.985 ;
  LAYER M1 ;
        RECT 14.925 19.235 15.175 20.245 ;
  LAYER M1 ;
        RECT 14.925 21.335 15.175 22.345 ;
  LAYER M1 ;
        RECT 14.495 15.455 14.745 18.985 ;
  LAYER M2 ;
        RECT 14.88 21.7 16.08 21.98 ;
  LAYER M2 ;
        RECT 15.74 15.4 16.94 15.68 ;
  LAYER M2 ;
        RECT 14.88 15.82 16.08 16.1 ;
  LAYER M2 ;
        RECT 15.74 19.6 16.94 19.88 ;
  LAYER M2 ;
        RECT 14.88 20.02 16.08 20.3 ;
  LAYER M2 ;
        RECT 14.45 16.24 16.51 16.52 ;
  LAYER M1 ;
        RECT 23.955 15.455 24.205 18.985 ;
  LAYER M1 ;
        RECT 23.955 19.235 24.205 20.245 ;
  LAYER M1 ;
        RECT 23.955 21.335 24.205 22.345 ;
  LAYER M1 ;
        RECT 17.935 15.455 18.185 18.985 ;
  LAYER M1 ;
        RECT 29.975 15.455 30.225 18.985 ;
  LAYER M2 ;
        RECT 17.89 15.4 30.27 15.68 ;
  LAYER M2 ;
        RECT 23.48 21.7 24.68 21.98 ;
  LAYER M2 ;
        RECT 23.48 15.82 24.68 16.1 ;
  LAYER M2 ;
        RECT 23.05 19.6 24.25 19.88 ;
  LAYER M3 ;
        RECT 24.37 15.38 24.65 22 ;
  LAYER M1 ;
        RECT 6.755 15.455 7.005 18.985 ;
  LAYER M1 ;
        RECT 6.755 19.235 7.005 20.245 ;
  LAYER M1 ;
        RECT 6.755 21.335 7.005 22.345 ;
  LAYER M1 ;
        RECT 12.775 15.455 13.025 18.985 ;
  LAYER M1 ;
        RECT 0.735 15.455 0.985 18.985 ;
  LAYER M2 ;
        RECT 0.69 15.4 13.07 15.68 ;
  LAYER M2 ;
        RECT 6.28 21.7 7.48 21.98 ;
  LAYER M2 ;
        RECT 6.28 15.82 7.48 16.1 ;
  LAYER M2 ;
        RECT 6.71 19.6 7.91 19.88 ;
  LAYER M3 ;
        RECT 6.31 15.38 6.59 22 ;
  END 
END DCDC_HUNIT_CONV2TO1
