MACRO CCP_PMOS_B_53083828_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CCP_PMOS_B_53083828_X1_Y1 0 0 ;
  SIZE 3440 BY 7560 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 6580 2320 6860 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1150 260 1430 4780 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 680 1860 5200 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 690 1120 2750 1400 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 7225 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M2 ;
      RECT 260 280 1460 560 ;
    LAYER M2 ;
      RECT 1120 4480 2320 4760 ;
    LAYER M2 ;
      RECT 1120 700 2320 980 ;
    LAYER M2 ;
      RECT 690 4900 1890 5180 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4955 1375 5125 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 2065 755 2235 925 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 1635 1175 1805 1345 ;
    LAYER V1 ;
      RECT 2495 1175 2665 1345 ;
    LAYER V2 ;
      RECT 1215 345 1365 495 ;
    LAYER V2 ;
      RECT 1215 4545 1365 4695 ;
    LAYER V2 ;
      RECT 1645 765 1795 915 ;
    LAYER V2 ;
      RECT 1645 4965 1795 5115 ;
    LAYER V0 ;
      RECT 1205 2705 1375 2875 ;
    LAYER V0 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V0 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V0 ;
      RECT 775 2705 945 2875 ;
    LAYER V0 ;
      RECT 1635 2705 1805 2875 ;
    LAYER V0 ;
      RECT 1635 2705 1805 2875 ;
    LAYER V0 ;
      RECT 2065 2705 2235 2875 ;
    LAYER V0 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V0 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V0 ;
      RECT 2495 2705 2665 2875 ;
  END
END CCP_PMOS_B_53083828_X1_Y1
MACRO DP_PMOS_B_25364157_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DP_PMOS_B_25364157_X1_Y1 0 0 ;
  SIZE 3440 BY 7560 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 6580 2320 6860 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260 280 1460 560 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 700 2320 980 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260 4480 1460 4760 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 4900 2320 5180 ;
    END
  END GB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 690 1120 2750 1400 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 7225 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 2065 755 2235 925 ;
    LAYER V1 ;
      RECT 2065 4955 2235 5125 ;
    LAYER V1 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 1635 1175 1805 1345 ;
    LAYER V1 ;
      RECT 2495 1175 2665 1345 ;
    LAYER V0 ;
      RECT 1205 2285 1375 2455 ;
    LAYER V0 ;
      RECT 1205 2625 1375 2795 ;
    LAYER V0 ;
      RECT 1205 2965 1375 3135 ;
    LAYER V0 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V0 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V0 ;
      RECT 775 2285 945 2455 ;
    LAYER V0 ;
      RECT 775 2625 945 2795 ;
    LAYER V0 ;
      RECT 775 2965 945 3135 ;
    LAYER V0 ;
      RECT 1635 2285 1805 2455 ;
    LAYER V0 ;
      RECT 1635 2285 1805 2455 ;
    LAYER V0 ;
      RECT 1635 2625 1805 2795 ;
    LAYER V0 ;
      RECT 1635 2625 1805 2795 ;
    LAYER V0 ;
      RECT 1635 2965 1805 3135 ;
    LAYER V0 ;
      RECT 1635 2965 1805 3135 ;
    LAYER V0 ;
      RECT 2065 2285 2235 2455 ;
    LAYER V0 ;
      RECT 2065 2625 2235 2795 ;
    LAYER V0 ;
      RECT 2065 2965 2235 3135 ;
    LAYER V0 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V0 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V0 ;
      RECT 2495 2285 2665 2455 ;
    LAYER V0 ;
      RECT 2495 2625 2665 2795 ;
    LAYER V0 ;
      RECT 2495 2965 2665 3135 ;
  END
END DP_PMOS_B_25364157_X1_Y1
MACRO DCAP_PMOS_57222488_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DCAP_PMOS_57222488_X1_Y1 0 0 ;
  SIZE 13760 BY 7560 ;
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5850 4480 7050 4760 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 7170 260 7450 6880 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 6755 4115 7005 5125 ;
    LAYER M1 ;
      RECT 6755 6215 7005 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 12775 335 13025 3865 ;
    LAYER M2 ;
      RECT 690 280 13070 560 ;
    LAYER M2 ;
      RECT 6280 6580 7480 6860 ;
    LAYER M2 ;
      RECT 6280 700 7480 980 ;
    LAYER V1 ;
      RECT 6795 755 6965 925 ;
    LAYER V1 ;
      RECT 6795 4535 6965 4705 ;
    LAYER V1 ;
      RECT 6795 6635 6965 6805 ;
    LAYER V1 ;
      RECT 775 335 945 505 ;
    LAYER V1 ;
      RECT 12815 335 12985 505 ;
    LAYER V2 ;
      RECT 7235 345 7385 495 ;
    LAYER V2 ;
      RECT 7235 765 7385 915 ;
    LAYER V2 ;
      RECT 7235 6645 7385 6795 ;
    LAYER V0 ;
      RECT 6795 1865 6965 2035 ;
    LAYER V0 ;
      RECT 6795 2205 6965 2375 ;
    LAYER V0 ;
      RECT 6795 2545 6965 2715 ;
    LAYER V0 ;
      RECT 6795 2885 6965 3055 ;
    LAYER V0 ;
      RECT 6795 3225 6965 3395 ;
    LAYER V0 ;
      RECT 6795 4535 6965 4705 ;
    LAYER V0 ;
      RECT 6795 6635 6965 6805 ;
    LAYER V0 ;
      RECT 775 1865 945 2035 ;
    LAYER V0 ;
      RECT 775 2205 945 2375 ;
    LAYER V0 ;
      RECT 775 2545 945 2715 ;
    LAYER V0 ;
      RECT 775 2885 945 3055 ;
    LAYER V0 ;
      RECT 775 3225 945 3395 ;
    LAYER V0 ;
      RECT 12815 1865 12985 2035 ;
    LAYER V0 ;
      RECT 12815 2205 12985 2375 ;
    LAYER V0 ;
      RECT 12815 2545 12985 2715 ;
    LAYER V0 ;
      RECT 12815 2885 12985 3055 ;
    LAYER V0 ;
      RECT 12815 3225 12985 3395 ;
  END
END DCAP_PMOS_57222488_X1_Y1
MACRO CCP_NMOS_B_26073270_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CCP_NMOS_B_26073270_X1_Y1 0 0 ;
  SIZE 3440 BY 7560 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 6580 2320 6860 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1150 260 1430 4780 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 680 1860 5200 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 690 1120 2750 1400 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 7225 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M2 ;
      RECT 260 280 1460 560 ;
    LAYER M2 ;
      RECT 1120 4480 2320 4760 ;
    LAYER M2 ;
      RECT 1120 700 2320 980 ;
    LAYER M2 ;
      RECT 690 4900 1890 5180 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4955 1375 5125 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 2065 755 2235 925 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 1635 1175 1805 1345 ;
    LAYER V1 ;
      RECT 2495 1175 2665 1345 ;
    LAYER V2 ;
      RECT 1215 345 1365 495 ;
    LAYER V2 ;
      RECT 1215 4545 1365 4695 ;
    LAYER V2 ;
      RECT 1645 765 1795 915 ;
    LAYER V2 ;
      RECT 1645 4965 1795 5115 ;
    LAYER V0 ;
      RECT 1205 2705 1375 2875 ;
    LAYER V0 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V0 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V0 ;
      RECT 775 2705 945 2875 ;
    LAYER V0 ;
      RECT 1635 2705 1805 2875 ;
    LAYER V0 ;
      RECT 1635 2705 1805 2875 ;
    LAYER V0 ;
      RECT 2065 2705 2235 2875 ;
    LAYER V0 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V0 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V0 ;
      RECT 2495 2705 2665 2875 ;
  END
END CCP_NMOS_B_26073270_X1_Y1
MACRO DP_NMOS_B_83449181_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_83449181_X1_Y1 0 0 ;
  SIZE 3440 BY 7560 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 6580 2320 6860 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260 280 1460 560 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 700 2320 980 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260 4480 1460 4760 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 4900 2320 5180 ;
    END
  END GB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 690 1120 2750 1400 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 7225 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 2065 755 2235 925 ;
    LAYER V1 ;
      RECT 2065 4955 2235 5125 ;
    LAYER V1 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 1635 1175 1805 1345 ;
    LAYER V1 ;
      RECT 2495 1175 2665 1345 ;
    LAYER V0 ;
      RECT 1205 2495 1375 2665 ;
    LAYER V0 ;
      RECT 1205 2835 1375 3005 ;
    LAYER V0 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V0 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V0 ;
      RECT 775 2495 945 2665 ;
    LAYER V0 ;
      RECT 775 2835 945 3005 ;
    LAYER V0 ;
      RECT 1635 2495 1805 2665 ;
    LAYER V0 ;
      RECT 1635 2495 1805 2665 ;
    LAYER V0 ;
      RECT 1635 2835 1805 3005 ;
    LAYER V0 ;
      RECT 1635 2835 1805 3005 ;
    LAYER V0 ;
      RECT 2065 2495 2235 2665 ;
    LAYER V0 ;
      RECT 2065 2835 2235 3005 ;
    LAYER V0 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V0 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V0 ;
      RECT 2495 2495 2665 2665 ;
    LAYER V0 ;
      RECT 2495 2835 2665 3005 ;
  END
END DP_NMOS_B_83449181_X1_Y1
