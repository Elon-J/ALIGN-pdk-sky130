MACRO PMOS_4T_43971774_X2_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN PMOS_4T_43971774_X2_Y1 0 0 ;
  SIZE 5160 BY 9240 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 7420 3180 7700 ;
    END
  END B
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 1120 3180 1400 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 5320 3180 5600 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1550 1540 3610 1820 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 2025 1175 2275 4705 ;
    LAYER M1 ;
      RECT 2025 4955 2275 5965 ;
    LAYER M1 ;
      RECT 2025 7055 2275 8065 ;
    LAYER M1 ;
      RECT 1595 1175 1845 4705 ;
    LAYER M1 ;
      RECT 2455 1175 2705 4705 ;
    LAYER M1 ;
      RECT 2885 1175 3135 4705 ;
    LAYER M1 ;
      RECT 2885 4955 3135 5965 ;
    LAYER M1 ;
      RECT 2885 7055 3135 8065 ;
    LAYER M1 ;
      RECT 3315 1175 3565 4705 ;
    LAYER V1 ;
      RECT 2065 1175 2235 1345 ;
    LAYER V1 ;
      RECT 2065 5375 2235 5545 ;
    LAYER V1 ;
      RECT 2065 7475 2235 7645 ;
    LAYER V1 ;
      RECT 2925 1175 3095 1345 ;
    LAYER V1 ;
      RECT 2925 5375 3095 5545 ;
    LAYER V1 ;
      RECT 2925 7475 3095 7645 ;
    LAYER V1 ;
      RECT 1635 1595 1805 1765 ;
    LAYER V1 ;
      RECT 2495 1595 2665 1765 ;
    LAYER V1 ;
      RECT 3355 1595 3525 1765 ;
    LAYER V0 ;
      RECT 2065 3545 2235 3715 ;
    LAYER V0 ;
      RECT 2065 5375 2235 5545 ;
    LAYER V0 ;
      RECT 2065 7475 2235 7645 ;
    LAYER V0 ;
      RECT 1635 3545 1805 3715 ;
    LAYER V0 ;
      RECT 2495 3545 2665 3715 ;
    LAYER V0 ;
      RECT 2495 3545 2665 3715 ;
    LAYER V0 ;
      RECT 2925 3545 3095 3715 ;
    LAYER V0 ;
      RECT 2925 5375 3095 5545 ;
    LAYER V0 ;
      RECT 2925 7475 3095 7645 ;
    LAYER V0 ;
      RECT 3355 3545 3525 3715 ;
  END
END PMOS_4T_43971774_X2_Y1
