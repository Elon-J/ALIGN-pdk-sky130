MACRO DCDC_DAC
  ORIGIN 0 0 ;
  FOREIGN DCDC_DAC 0 0 ;
  SIZE 14.62 BY 22.68 ;
  PIN D0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
      LAYER M2 ;
        RECT 6.28 2.8 7.48 3.08 ;
      LAYER M2 ;
        RECT 4.73 2.8 6.45 3.08 ;
    END
  END D0
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 6.28 0.7 7.48 0.98 ;
      LAYER M2 ;
        RECT 6.28 15.82 7.48 16.1 ;
      LAYER M2 ;
        RECT 9.72 0.7 10.92 0.98 ;
      LAYER M2 ;
        RECT 6.28 8.26 7.48 8.54 ;
      LAYER M2 ;
        RECT 9.72 8.26 10.92 8.54 ;
      LAYER M2 ;
        RECT 9.72 15.82 10.92 16.1 ;
      LAYER M2 ;
        RECT 6.72 0.7 7.04 0.98 ;
      LAYER M3 ;
        RECT 6.74 0.84 7.02 15.96 ;
      LAYER M2 ;
        RECT 6.72 15.82 7.04 16.1 ;
      LAYER M2 ;
        RECT 7.31 0.7 9.89 0.98 ;
      LAYER M3 ;
        RECT 6.74 8.215 7.02 8.585 ;
      LAYER M2 ;
        RECT 6.72 8.26 7.04 8.54 ;
      LAYER M2 ;
        RECT 7.31 8.26 9.89 8.54 ;
      LAYER M2 ;
        RECT 7.31 15.82 9.89 16.1 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
      LAYER M3 ;
        RECT 3.3 15.8 3.58 22 ;
      LAYER M3 ;
        RECT 13.62 0.68 13.9 6.88 ;
      LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
      LAYER M3 ;
        RECT 13.62 8.24 13.9 14.44 ;
      LAYER M3 ;
        RECT 13.62 15.8 13.9 22 ;
      LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
      LAYER M3 ;
        RECT 3.3 6.72 3.58 7.56 ;
      LAYER M2 ;
        RECT 3.01 7.42 3.44 7.7 ;
      LAYER M1 ;
        RECT 2.885 7.56 3.135 15.12 ;
      LAYER M2 ;
        RECT 3.01 14.98 3.44 15.26 ;
      LAYER M3 ;
        RECT 3.3 15.12 3.58 15.96 ;
      LAYER M3 ;
        RECT 3.3 3.595 3.58 3.965 ;
      LAYER M2 ;
        RECT 3.44 3.64 13.76 3.92 ;
      LAYER M3 ;
        RECT 13.62 3.595 13.9 3.965 ;
      LAYER M1 ;
        RECT 2.885 11.255 3.135 11.425 ;
      LAYER M2 ;
        RECT 3.01 11.2 3.44 11.48 ;
      LAYER M3 ;
        RECT 3.3 11.155 3.58 11.525 ;
      LAYER M3 ;
        RECT 13.62 6.72 13.9 8.4 ;
      LAYER M3 ;
        RECT 13.62 14.28 13.9 15.96 ;
      LAYER M3 ;
        RECT 3.3 3.595 3.58 3.965 ;
      LAYER M4 ;
        RECT 1.72 3.38 3.44 4.18 ;
      LAYER M3 ;
        RECT 1.58 3.595 1.86 3.965 ;
    END
  END VGND
  PIN REF
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 5.85 6.58 7.91 6.86 ;
      LAYER M2 ;
        RECT 5.85 21.7 7.91 21.98 ;
      LAYER M2 ;
        RECT 9.29 6.58 11.35 6.86 ;
      LAYER M2 ;
        RECT 5.85 14.14 7.91 14.42 ;
      LAYER M2 ;
        RECT 9.29 14.14 11.35 14.42 ;
      LAYER M2 ;
        RECT 9.29 21.7 11.35 21.98 ;
      LAYER M2 ;
        RECT 6.29 6.58 6.61 6.86 ;
      LAYER M3 ;
        RECT 6.31 6.72 6.59 21.84 ;
      LAYER M2 ;
        RECT 6.29 21.7 6.61 21.98 ;
      LAYER M2 ;
        RECT 7.74 6.58 9.46 6.86 ;
      LAYER M3 ;
        RECT 6.31 14.095 6.59 14.465 ;
      LAYER M2 ;
        RECT 6.29 14.14 6.61 14.42 ;
      LAYER M2 ;
        RECT 7.74 14.14 9.46 14.42 ;
      LAYER M2 ;
        RECT 7.74 21.7 9.46 21.98 ;
    END
  END REF
  PIN D5
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.7 17.92 4.9 18.2 ;
      LAYER M2 ;
        RECT 6.28 17.92 7.48 18.2 ;
      LAYER M2 ;
        RECT 4.73 17.92 6.45 18.2 ;
    END
  END D5
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 12.3 2.8 13.5 3.08 ;
      LAYER M2 ;
        RECT 9.72 2.8 10.92 3.08 ;
      LAYER M2 ;
        RECT 10.75 2.8 12.47 3.08 ;
    END
  END D1
  PIN D2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.7 10.36 4.9 10.64 ;
      LAYER M2 ;
        RECT 6.28 10.36 7.48 10.64 ;
      LAYER M2 ;
        RECT 4.73 10.36 6.45 10.64 ;
    END
  END D2
  PIN D3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 12.3 10.36 13.5 10.64 ;
      LAYER M2 ;
        RECT 9.72 10.36 10.92 10.64 ;
      LAYER M2 ;
        RECT 10.75 10.36 12.47 10.64 ;
    END
  END D3
  PIN D4
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 12.3 17.92 13.5 18.2 ;
      LAYER M2 ;
        RECT 9.72 17.92 10.92 18.2 ;
      LAYER M2 ;
        RECT 10.75 17.92 12.47 18.2 ;
    END
  END D4
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.26 0.28 1.46 0.56 ;
    END
  END VOUT
  PIN RST
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.26 4.48 1.46 4.76 ;
    END
  END RST
  OBS 
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 6.28 7 7.48 7.28 ;
  LAYER M2 ;
        RECT 4.73 7 6.45 7.28 ;
  LAYER M2 ;
        RECT 3.7 22.12 4.9 22.4 ;
  LAYER M2 ;
        RECT 6.28 22.12 7.48 22.4 ;
  LAYER M2 ;
        RECT 4.73 22.12 6.45 22.4 ;
  LAYER M2 ;
        RECT 12.3 7 13.5 7.28 ;
  LAYER M2 ;
        RECT 9.72 7 10.92 7.28 ;
  LAYER M2 ;
        RECT 10.75 7 12.47 7.28 ;
  LAYER M2 ;
        RECT 3.7 14.56 4.9 14.84 ;
  LAYER M2 ;
        RECT 6.28 14.56 7.48 14.84 ;
  LAYER M2 ;
        RECT 4.73 14.56 6.45 14.84 ;
  LAYER M2 ;
        RECT 12.3 14.56 13.5 14.84 ;
  LAYER M2 ;
        RECT 9.72 14.56 10.92 14.84 ;
  LAYER M2 ;
        RECT 10.75 14.56 12.47 14.84 ;
  LAYER M2 ;
        RECT 12.3 22.12 13.5 22.4 ;
  LAYER M2 ;
        RECT 9.72 22.12 10.92 22.4 ;
  LAYER M2 ;
        RECT 10.75 22.12 12.47 22.4 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M2 ;
        RECT 3.27 6.58 4.47 6.86 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
  LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M2 ;
        RECT 6.28 0.7 7.48 0.98 ;
  LAYER M2 ;
        RECT 6.28 7 7.48 7.28 ;
  LAYER M2 ;
        RECT 6.28 2.8 7.48 3.08 ;
  LAYER M2 ;
        RECT 5.85 6.58 7.91 6.86 ;
  LAYER M1 ;
        RECT 3.745 18.815 3.995 22.345 ;
  LAYER M1 ;
        RECT 3.745 17.555 3.995 18.565 ;
  LAYER M1 ;
        RECT 3.745 15.455 3.995 16.465 ;
  LAYER M1 ;
        RECT 4.175 18.815 4.425 22.345 ;
  LAYER M1 ;
        RECT 3.315 18.815 3.565 22.345 ;
  LAYER M2 ;
        RECT 3.27 21.7 4.47 21.98 ;
  LAYER M2 ;
        RECT 3.27 15.82 4.47 16.1 ;
  LAYER M2 ;
        RECT 3.7 22.12 4.9 22.4 ;
  LAYER M2 ;
        RECT 3.7 17.92 4.9 18.2 ;
  LAYER M3 ;
        RECT 3.3 15.8 3.58 22 ;
  LAYER M1 ;
        RECT 7.185 18.815 7.435 22.345 ;
  LAYER M1 ;
        RECT 7.185 17.555 7.435 18.565 ;
  LAYER M1 ;
        RECT 7.185 15.455 7.435 16.465 ;
  LAYER M1 ;
        RECT 7.615 18.815 7.865 22.345 ;
  LAYER M1 ;
        RECT 6.755 18.815 7.005 22.345 ;
  LAYER M1 ;
        RECT 6.325 18.815 6.575 22.345 ;
  LAYER M1 ;
        RECT 6.325 17.555 6.575 18.565 ;
  LAYER M1 ;
        RECT 6.325 15.455 6.575 16.465 ;
  LAYER M1 ;
        RECT 5.895 18.815 6.145 22.345 ;
  LAYER M2 ;
        RECT 6.28 15.82 7.48 16.1 ;
  LAYER M2 ;
        RECT 6.28 22.12 7.48 22.4 ;
  LAYER M2 ;
        RECT 6.28 17.92 7.48 18.2 ;
  LAYER M2 ;
        RECT 5.85 21.7 7.91 21.98 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M2 ;
        RECT 12.73 6.58 13.93 6.86 ;
  LAYER M2 ;
        RECT 12.73 0.7 13.93 0.98 ;
  LAYER M2 ;
        RECT 12.3 7 13.5 7.28 ;
  LAYER M2 ;
        RECT 12.3 2.8 13.5 3.08 ;
  LAYER M3 ;
        RECT 13.62 0.68 13.9 6.88 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 10.625 2.435 10.875 3.445 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 1.345 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M2 ;
        RECT 9.72 0.7 10.92 0.98 ;
  LAYER M2 ;
        RECT 9.72 7 10.92 7.28 ;
  LAYER M2 ;
        RECT 9.72 2.8 10.92 3.08 ;
  LAYER M2 ;
        RECT 9.29 6.58 11.35 6.86 ;
  LAYER M1 ;
        RECT 3.745 11.255 3.995 14.785 ;
  LAYER M1 ;
        RECT 3.745 9.995 3.995 11.005 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 8.905 ;
  LAYER M1 ;
        RECT 4.175 11.255 4.425 14.785 ;
  LAYER M1 ;
        RECT 3.315 11.255 3.565 14.785 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 3.7 14.56 4.9 14.84 ;
  LAYER M2 ;
        RECT 3.7 10.36 4.9 10.64 ;
  LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
  LAYER M1 ;
        RECT 7.185 11.255 7.435 14.785 ;
  LAYER M1 ;
        RECT 7.185 9.995 7.435 11.005 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 8.905 ;
  LAYER M1 ;
        RECT 7.615 11.255 7.865 14.785 ;
  LAYER M1 ;
        RECT 6.755 11.255 7.005 14.785 ;
  LAYER M1 ;
        RECT 6.325 11.255 6.575 14.785 ;
  LAYER M1 ;
        RECT 6.325 9.995 6.575 11.005 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 8.905 ;
  LAYER M1 ;
        RECT 5.895 11.255 6.145 14.785 ;
  LAYER M2 ;
        RECT 6.28 8.26 7.48 8.54 ;
  LAYER M2 ;
        RECT 6.28 14.56 7.48 14.84 ;
  LAYER M2 ;
        RECT 6.28 10.36 7.48 10.64 ;
  LAYER M2 ;
        RECT 5.85 14.14 7.91 14.42 ;
  LAYER M1 ;
        RECT 13.205 11.255 13.455 14.785 ;
  LAYER M1 ;
        RECT 13.205 9.995 13.455 11.005 ;
  LAYER M1 ;
        RECT 13.205 7.895 13.455 8.905 ;
  LAYER M1 ;
        RECT 12.775 11.255 13.025 14.785 ;
  LAYER M1 ;
        RECT 13.635 11.255 13.885 14.785 ;
  LAYER M2 ;
        RECT 12.73 14.14 13.93 14.42 ;
  LAYER M2 ;
        RECT 12.73 8.26 13.93 8.54 ;
  LAYER M2 ;
        RECT 12.3 14.56 13.5 14.84 ;
  LAYER M2 ;
        RECT 12.3 10.36 13.5 10.64 ;
  LAYER M3 ;
        RECT 13.62 8.24 13.9 14.44 ;
  LAYER M1 ;
        RECT 9.765 11.255 10.015 14.785 ;
  LAYER M1 ;
        RECT 9.765 9.995 10.015 11.005 ;
  LAYER M1 ;
        RECT 9.765 7.895 10.015 8.905 ;
  LAYER M1 ;
        RECT 9.335 11.255 9.585 14.785 ;
  LAYER M1 ;
        RECT 10.195 11.255 10.445 14.785 ;
  LAYER M1 ;
        RECT 10.625 11.255 10.875 14.785 ;
  LAYER M1 ;
        RECT 10.625 9.995 10.875 11.005 ;
  LAYER M1 ;
        RECT 10.625 7.895 10.875 8.905 ;
  LAYER M1 ;
        RECT 11.055 11.255 11.305 14.785 ;
  LAYER M2 ;
        RECT 9.72 8.26 10.92 8.54 ;
  LAYER M2 ;
        RECT 9.72 14.56 10.92 14.84 ;
  LAYER M2 ;
        RECT 9.72 10.36 10.92 10.64 ;
  LAYER M2 ;
        RECT 9.29 14.14 11.35 14.42 ;
  LAYER M1 ;
        RECT 13.205 18.815 13.455 22.345 ;
  LAYER M1 ;
        RECT 13.205 17.555 13.455 18.565 ;
  LAYER M1 ;
        RECT 13.205 15.455 13.455 16.465 ;
  LAYER M1 ;
        RECT 12.775 18.815 13.025 22.345 ;
  LAYER M1 ;
        RECT 13.635 18.815 13.885 22.345 ;
  LAYER M2 ;
        RECT 12.73 21.7 13.93 21.98 ;
  LAYER M2 ;
        RECT 12.73 15.82 13.93 16.1 ;
  LAYER M2 ;
        RECT 12.3 22.12 13.5 22.4 ;
  LAYER M2 ;
        RECT 12.3 17.92 13.5 18.2 ;
  LAYER M3 ;
        RECT 13.62 15.8 13.9 22 ;
  LAYER M1 ;
        RECT 9.765 18.815 10.015 22.345 ;
  LAYER M1 ;
        RECT 9.765 17.555 10.015 18.565 ;
  LAYER M1 ;
        RECT 9.765 15.455 10.015 16.465 ;
  LAYER M1 ;
        RECT 9.335 18.815 9.585 22.345 ;
  LAYER M1 ;
        RECT 10.195 18.815 10.445 22.345 ;
  LAYER M1 ;
        RECT 10.625 18.815 10.875 22.345 ;
  LAYER M1 ;
        RECT 10.625 17.555 10.875 18.565 ;
  LAYER M1 ;
        RECT 10.625 15.455 10.875 16.465 ;
  LAYER M1 ;
        RECT 11.055 18.815 11.305 22.345 ;
  LAYER M2 ;
        RECT 9.72 15.82 10.92 16.1 ;
  LAYER M2 ;
        RECT 9.72 22.12 10.92 22.4 ;
  LAYER M2 ;
        RECT 9.72 17.92 10.92 18.2 ;
  LAYER M2 ;
        RECT 9.29 21.7 11.35 21.98 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 3.865 ;
  LAYER M1 ;
        RECT 1.165 4.115 1.415 5.125 ;
  LAYER M1 ;
        RECT 1.165 6.215 1.415 7.225 ;
  LAYER M1 ;
        RECT 0.735 0.335 0.985 3.865 ;
  LAYER M1 ;
        RECT 1.595 0.335 1.845 3.865 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 0.69 6.58 1.89 6.86 ;
  LAYER M2 ;
        RECT 0.26 0.28 1.46 0.56 ;
  LAYER M2 ;
        RECT 0.26 4.48 1.46 4.76 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
  END 
END DCDC_DAC
