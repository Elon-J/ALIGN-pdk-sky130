MACRO DCDC_CONV2TO1_1
  ORIGIN 0 0 ;
  FOREIGN DCDC_CONV2TO1_1 0 0 ;
  SIZE 64.07 BY 31.5 ;
  PIN CLK0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 6.31 16.22 6.59 22.84 ;
      LAYER M3 ;
        RECT 57.48 16.22 57.76 22.84 ;
      LAYER M3 ;
        RECT 6.31 16.195 6.59 16.565 ;
      LAYER M4 ;
        RECT 6.45 15.98 57.62 16.78 ;
      LAYER M3 ;
        RECT 57.48 16.195 57.76 16.565 ;
    END
  END CLK0
  PIN CLK0B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 25.23 8.66 25.51 15.28 ;
      LAYER M3 ;
        RECT 38.56 8.66 38.84 15.28 ;
      LAYER M3 ;
        RECT 25.23 11.155 25.51 11.525 ;
      LAYER M4 ;
        RECT 25.37 10.94 38.7 11.74 ;
      LAYER M3 ;
        RECT 38.56 11.155 38.84 11.525 ;
    END
  END CLK0B
  PIN CLK1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 25.23 16.22 25.51 22.84 ;
      LAYER M3 ;
        RECT 38.56 16.22 38.84 22.84 ;
      LAYER M3 ;
        RECT 25.23 15.96 25.51 16.38 ;
      LAYER M2 ;
        RECT 25.37 15.82 25.8 16.1 ;
      LAYER M3 ;
        RECT 25.66 15.12 25.94 15.96 ;
      LAYER M4 ;
        RECT 25.8 14.72 34.4 15.52 ;
      LAYER M3 ;
        RECT 34.26 15.12 34.54 15.96 ;
      LAYER M2 ;
        RECT 34.4 15.82 38.7 16.1 ;
      LAYER M3 ;
        RECT 38.56 15.96 38.84 16.38 ;
    END
  END CLK1
  PIN CLK1B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 6.31 8.66 6.59 15.28 ;
      LAYER M3 ;
        RECT 57.48 8.66 57.76 15.28 ;
      LAYER M3 ;
        RECT 6.31 14.935 6.59 15.305 ;
      LAYER M4 ;
        RECT 6.45 14.72 6.88 15.52 ;
      LAYER M3 ;
        RECT 6.74 15.12 7.02 17.64 ;
      LAYER M4 ;
        RECT 6.88 17.24 51.6 18.04 ;
      LAYER M3 ;
        RECT 51.46 15.54 51.74 17.64 ;
      LAYER M2 ;
        RECT 51.6 15.4 57.62 15.68 ;
      LAYER M3 ;
        RECT 57.48 15.12 57.76 15.54 ;
    END
  END CLK1B
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.31 30.52 16.51 30.8 ;
      LAYER M2 ;
        RECT 15.31 22.54 16.51 22.82 ;
      LAYER M2 ;
        RECT 15.32 30.52 15.64 30.8 ;
      LAYER M3 ;
        RECT 15.34 22.68 15.62 30.66 ;
      LAYER M2 ;
        RECT 15.32 22.54 15.64 22.82 ;
      LAYER M2 ;
        RECT 47.56 30.52 48.76 30.8 ;
      LAYER M2 ;
        RECT 47.56 22.54 48.76 22.82 ;
      LAYER M2 ;
        RECT 48.43 30.52 48.75 30.8 ;
      LAYER M3 ;
        RECT 48.45 22.68 48.73 30.66 ;
      LAYER M2 ;
        RECT 48.43 22.54 48.75 22.82 ;
      LAYER M2 ;
        RECT 16.34 22.54 16.77 22.82 ;
      LAYER M3 ;
        RECT 16.63 22.559 16.91 22.801 ;
      LAYER M4 ;
        RECT 16.77 22.28 43 23.08 ;
      LAYER M3 ;
        RECT 42.86 22.559 43.14 22.801 ;
      LAYER M2 ;
        RECT 43 22.54 47.73 22.82 ;
    END
  END VGND
  PIN VHIGH
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.88 6.16 16.94 6.44 ;
      LAYER M2 ;
        RECT 14.88 14.14 16.94 14.42 ;
      LAYER M2 ;
        RECT 14.89 6.16 15.21 6.44 ;
      LAYER M3 ;
        RECT 14.91 6.3 15.19 14.28 ;
      LAYER M2 ;
        RECT 14.89 14.14 15.21 14.42 ;
    END
  END VHIGH
  PIN VMID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.88 25.06 16.94 25.34 ;
      LAYER M2 ;
        RECT 14.88 17.08 16.94 17.36 ;
      LAYER M2 ;
        RECT 14.89 25.06 15.21 25.34 ;
      LAYER M3 ;
        RECT 14.91 17.22 15.19 25.2 ;
      LAYER M2 ;
        RECT 14.89 17.08 15.21 17.36 ;
      LAYER M2 ;
        RECT 47.13 6.16 49.19 6.44 ;
      LAYER M2 ;
        RECT 47.13 14.14 49.19 14.42 ;
      LAYER M2 ;
        RECT 48.86 6.16 49.18 6.44 ;
      LAYER M3 ;
        RECT 48.88 6.3 49.16 14.28 ;
      LAYER M2 ;
        RECT 48.86 14.14 49.18 14.42 ;
      LAYER M2 ;
        RECT 16.77 17.08 17.2 17.36 ;
      LAYER M3 ;
        RECT 17.06 15.54 17.34 17.22 ;
      LAYER M2 ;
        RECT 17.2 15.4 43 15.68 ;
      LAYER M1 ;
        RECT 42.875 14.28 43.125 15.54 ;
      LAYER M2 ;
        RECT 43 14.14 47.3 14.42 ;
    END
  END VMID
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.31 0.7 16.51 0.98 ;
      LAYER M2 ;
        RECT 15.31 8.68 16.51 8.96 ;
      LAYER M2 ;
        RECT 15.32 0.7 15.64 0.98 ;
      LAYER M3 ;
        RECT 15.34 0.84 15.62 8.82 ;
      LAYER M2 ;
        RECT 15.32 8.68 15.64 8.96 ;
      LAYER M2 ;
        RECT 47.56 0.7 48.76 0.98 ;
      LAYER M2 ;
        RECT 47.56 8.68 48.76 8.96 ;
      LAYER M2 ;
        RECT 48.43 0.7 48.75 0.98 ;
      LAYER M3 ;
        RECT 48.45 0.84 48.73 8.82 ;
      LAYER M2 ;
        RECT 48.43 8.68 48.75 8.96 ;
      LAYER M2 ;
        RECT 16.34 8.68 16.77 8.96 ;
      LAYER M1 ;
        RECT 16.645 8.82 16.895 9.24 ;
      LAYER M2 ;
        RECT 16.77 9.1 43 9.38 ;
      LAYER M1 ;
        RECT 42.875 8.82 43.125 9.24 ;
      LAYER M2 ;
        RECT 43 8.68 47.73 8.96 ;
    END
  END VPWR
  PIN Y0_TOP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 16.17 14.98 17.37 15.26 ;
      LAYER M2 ;
        RECT 16.17 16.24 17.37 16.52 ;
      LAYER M2 ;
        RECT 16.61 14.98 16.93 15.26 ;
      LAYER M3 ;
        RECT 16.63 15.12 16.91 16.38 ;
      LAYER M2 ;
        RECT 16.61 16.24 16.93 16.52 ;
    END
  END Y0_TOP
  PIN Y1_TOP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.31 14.56 16.51 14.84 ;
      LAYER M2 ;
        RECT 15.31 16.66 16.51 16.94 ;
      LAYER M2 ;
        RECT 15.75 14.56 16.07 14.84 ;
      LAYER M3 ;
        RECT 15.77 14.7 16.05 16.8 ;
      LAYER M2 ;
        RECT 15.75 16.66 16.07 16.94 ;
    END
  END Y1_TOP
  PIN VLOW
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 47.13 25.06 49.19 25.34 ;
      LAYER M2 ;
        RECT 47.13 17.08 49.19 17.36 ;
      LAYER M2 ;
        RECT 48.86 25.06 49.18 25.34 ;
      LAYER M3 ;
        RECT 48.88 17.22 49.16 25.2 ;
      LAYER M2 ;
        RECT 48.86 17.08 49.18 17.36 ;
    END
  END VLOW
  PIN Y0_BOT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 46.7 14.98 47.9 15.26 ;
      LAYER M2 ;
        RECT 46.7 16.24 47.9 16.52 ;
      LAYER M2 ;
        RECT 47.14 14.98 47.46 15.26 ;
      LAYER M3 ;
        RECT 47.16 15.12 47.44 16.38 ;
      LAYER M2 ;
        RECT 47.14 16.24 47.46 16.52 ;
    END
  END Y0_BOT
  PIN Y1_BOT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 47.56 14.56 48.76 14.84 ;
      LAYER M2 ;
        RECT 47.56 16.66 48.76 16.94 ;
      LAYER M2 ;
        RECT 48 14.56 48.32 14.84 ;
      LAYER M3 ;
        RECT 48.02 14.7 48.3 16.8 ;
      LAYER M2 ;
        RECT 48 16.66 48.32 16.94 ;
    END
  END Y1_BOT
  OBS 
  LAYER M3 ;
        RECT 16.2 2.78 16.48 7.3 ;
  LAYER M2 ;
        RECT 16.17 10.78 17.37 11.06 ;
  LAYER M2 ;
        RECT 23.91 10.78 25.11 11.06 ;
  LAYER M3 ;
        RECT 16.2 7.14 16.48 10.92 ;
  LAYER M2 ;
        RECT 16.18 10.78 16.5 11.06 ;
  LAYER M2 ;
        RECT 17.2 10.78 24.08 11.06 ;
  LAYER M2 ;
        RECT 16.18 10.78 16.5 11.06 ;
  LAYER M3 ;
        RECT 16.2 10.76 16.48 11.08 ;
  LAYER M2 ;
        RECT 16.18 10.78 16.5 11.06 ;
  LAYER M3 ;
        RECT 16.2 10.76 16.48 11.08 ;
  LAYER M2 ;
        RECT 16.18 10.78 16.5 11.06 ;
  LAYER M3 ;
        RECT 16.2 10.76 16.48 11.08 ;
  LAYER M2 ;
        RECT 16.18 10.78 16.5 11.06 ;
  LAYER M3 ;
        RECT 16.2 10.76 16.48 11.08 ;
  LAYER M3 ;
        RECT 15.77 2.36 16.05 6.88 ;
  LAYER M2 ;
        RECT 15.31 10.36 16.51 10.64 ;
  LAYER M2 ;
        RECT 6.71 10.78 7.91 11.06 ;
  LAYER M3 ;
        RECT 15.77 6.72 16.05 10.5 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M2 ;
        RECT 15.32 10.36 15.64 10.64 ;
  LAYER M3 ;
        RECT 15.34 10.5 15.62 10.92 ;
  LAYER M2 ;
        RECT 7.74 10.78 15.48 11.06 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M2 ;
        RECT 15.32 10.36 15.64 10.64 ;
  LAYER M3 ;
        RECT 15.34 10.34 15.62 10.66 ;
  LAYER M2 ;
        RECT 15.32 10.78 15.64 11.06 ;
  LAYER M3 ;
        RECT 15.34 10.76 15.62 11.08 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M2 ;
        RECT 15.32 10.36 15.64 10.64 ;
  LAYER M3 ;
        RECT 15.34 10.34 15.62 10.66 ;
  LAYER M2 ;
        RECT 15.32 10.78 15.64 11.06 ;
  LAYER M3 ;
        RECT 15.34 10.76 15.62 11.08 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 16.215 2.435 16.465 3.445 ;
  LAYER M1 ;
        RECT 16.215 0.335 16.465 1.345 ;
  LAYER M1 ;
        RECT 16.645 3.695 16.895 7.225 ;
  LAYER M1 ;
        RECT 15.785 3.695 16.035 7.225 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M1 ;
        RECT 15.355 2.435 15.605 3.445 ;
  LAYER M1 ;
        RECT 15.355 0.335 15.605 1.345 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M2 ;
        RECT 16.17 7 17.37 7.28 ;
  LAYER M2 ;
        RECT 15.31 2.8 16.51 3.08 ;
  LAYER M2 ;
        RECT 15.31 6.58 16.51 6.86 ;
  LAYER M2 ;
        RECT 15.74 2.38 16.94 2.66 ;
  LAYER M2 ;
        RECT 15.31 0.7 16.51 0.98 ;
  LAYER M3 ;
        RECT 16.2 2.78 16.48 7.3 ;
  LAYER M3 ;
        RECT 15.77 2.36 16.05 6.88 ;
  LAYER M2 ;
        RECT 14.88 6.16 16.94 6.44 ;
  LAYER M1 ;
        RECT 16.215 11.675 16.465 15.205 ;
  LAYER M1 ;
        RECT 16.215 10.415 16.465 11.425 ;
  LAYER M1 ;
        RECT 16.215 8.315 16.465 9.325 ;
  LAYER M1 ;
        RECT 16.645 11.675 16.895 15.205 ;
  LAYER M1 ;
        RECT 15.785 11.675 16.035 15.205 ;
  LAYER M1 ;
        RECT 15.355 11.675 15.605 15.205 ;
  LAYER M1 ;
        RECT 15.355 10.415 15.605 11.425 ;
  LAYER M1 ;
        RECT 15.355 8.315 15.605 9.325 ;
  LAYER M1 ;
        RECT 14.925 11.675 15.175 15.205 ;
  LAYER M2 ;
        RECT 15.31 8.68 16.51 8.96 ;
  LAYER M2 ;
        RECT 16.17 14.98 17.37 15.26 ;
  LAYER M2 ;
        RECT 15.31 14.56 16.51 14.84 ;
  LAYER M2 ;
        RECT 16.17 10.78 17.37 11.06 ;
  LAYER M2 ;
        RECT 15.31 10.36 16.51 10.64 ;
  LAYER M2 ;
        RECT 14.88 14.14 16.94 14.42 ;
  LAYER M1 ;
        RECT 24.815 11.675 25.065 15.205 ;
  LAYER M1 ;
        RECT 24.815 10.415 25.065 11.425 ;
  LAYER M1 ;
        RECT 24.815 8.315 25.065 9.325 ;
  LAYER M1 ;
        RECT 18.795 11.675 19.045 15.205 ;
  LAYER M1 ;
        RECT 30.835 11.675 31.085 15.205 ;
  LAYER M2 ;
        RECT 24.34 14.98 25.54 15.26 ;
  LAYER M2 ;
        RECT 18.75 14.56 31.13 14.84 ;
  LAYER M2 ;
        RECT 24.34 8.68 25.54 8.96 ;
  LAYER M2 ;
        RECT 23.91 10.78 25.11 11.06 ;
  LAYER M3 ;
        RECT 25.23 8.66 25.51 15.28 ;
  LAYER M1 ;
        RECT 6.755 11.675 7.005 15.205 ;
  LAYER M1 ;
        RECT 6.755 10.415 7.005 11.425 ;
  LAYER M1 ;
        RECT 6.755 8.315 7.005 9.325 ;
  LAYER M1 ;
        RECT 12.775 11.675 13.025 15.205 ;
  LAYER M1 ;
        RECT 0.735 11.675 0.985 15.205 ;
  LAYER M2 ;
        RECT 6.28 14.98 7.48 15.26 ;
  LAYER M2 ;
        RECT 0.69 14.56 13.07 14.84 ;
  LAYER M2 ;
        RECT 6.28 8.68 7.48 8.96 ;
  LAYER M2 ;
        RECT 6.71 10.78 7.91 11.06 ;
  LAYER M3 ;
        RECT 6.31 8.66 6.59 15.28 ;
  LAYER M3 ;
        RECT 16.2 24.2 16.48 28.72 ;
  LAYER M2 ;
        RECT 16.17 20.44 17.37 20.72 ;
  LAYER M2 ;
        RECT 23.91 20.44 25.11 20.72 ;
  LAYER M3 ;
        RECT 16.2 20.58 16.48 24.36 ;
  LAYER M2 ;
        RECT 16.18 20.44 16.5 20.72 ;
  LAYER M2 ;
        RECT 17.2 20.44 24.08 20.72 ;
  LAYER M2 ;
        RECT 16.18 20.44 16.5 20.72 ;
  LAYER M3 ;
        RECT 16.2 20.42 16.48 20.74 ;
  LAYER M2 ;
        RECT 16.18 20.44 16.5 20.72 ;
  LAYER M3 ;
        RECT 16.2 20.42 16.48 20.74 ;
  LAYER M2 ;
        RECT 16.18 20.44 16.5 20.72 ;
  LAYER M3 ;
        RECT 16.2 20.42 16.48 20.74 ;
  LAYER M2 ;
        RECT 16.18 20.44 16.5 20.72 ;
  LAYER M3 ;
        RECT 16.2 20.42 16.48 20.74 ;
  LAYER M3 ;
        RECT 15.77 24.62 16.05 29.14 ;
  LAYER M2 ;
        RECT 15.31 20.86 16.51 21.14 ;
  LAYER M2 ;
        RECT 6.71 20.44 7.91 20.72 ;
  LAYER M3 ;
        RECT 15.77 21 16.05 24.78 ;
  LAYER M2 ;
        RECT 15.75 20.86 16.07 21.14 ;
  LAYER M2 ;
        RECT 15.32 20.86 15.64 21.14 ;
  LAYER M3 ;
        RECT 15.34 20.58 15.62 21 ;
  LAYER M2 ;
        RECT 7.74 20.44 15.48 20.72 ;
  LAYER M2 ;
        RECT 15.75 20.86 16.07 21.14 ;
  LAYER M3 ;
        RECT 15.77 20.84 16.05 21.16 ;
  LAYER M2 ;
        RECT 15.75 20.86 16.07 21.14 ;
  LAYER M3 ;
        RECT 15.77 20.84 16.05 21.16 ;
  LAYER M2 ;
        RECT 15.32 20.86 15.64 21.14 ;
  LAYER M3 ;
        RECT 15.34 20.84 15.62 21.16 ;
  LAYER M2 ;
        RECT 15.32 20.44 15.64 20.72 ;
  LAYER M3 ;
        RECT 15.34 20.42 15.62 20.74 ;
  LAYER M2 ;
        RECT 15.75 20.86 16.07 21.14 ;
  LAYER M3 ;
        RECT 15.77 20.84 16.05 21.16 ;
  LAYER M2 ;
        RECT 15.32 20.86 15.64 21.14 ;
  LAYER M3 ;
        RECT 15.34 20.84 15.62 21.16 ;
  LAYER M2 ;
        RECT 15.32 20.44 15.64 20.72 ;
  LAYER M3 ;
        RECT 15.34 20.42 15.62 20.74 ;
  LAYER M2 ;
        RECT 15.75 20.86 16.07 21.14 ;
  LAYER M3 ;
        RECT 15.77 20.84 16.05 21.16 ;
  LAYER M1 ;
        RECT 16.215 24.275 16.465 27.805 ;
  LAYER M1 ;
        RECT 16.215 28.055 16.465 29.065 ;
  LAYER M1 ;
        RECT 16.215 30.155 16.465 31.165 ;
  LAYER M1 ;
        RECT 16.645 24.275 16.895 27.805 ;
  LAYER M1 ;
        RECT 15.785 24.275 16.035 27.805 ;
  LAYER M1 ;
        RECT 15.355 24.275 15.605 27.805 ;
  LAYER M1 ;
        RECT 15.355 28.055 15.605 29.065 ;
  LAYER M1 ;
        RECT 15.355 30.155 15.605 31.165 ;
  LAYER M1 ;
        RECT 14.925 24.275 15.175 27.805 ;
  LAYER M2 ;
        RECT 16.17 24.22 17.37 24.5 ;
  LAYER M2 ;
        RECT 15.31 28.42 16.51 28.7 ;
  LAYER M2 ;
        RECT 15.31 24.64 16.51 24.92 ;
  LAYER M2 ;
        RECT 15.74 28.84 16.94 29.12 ;
  LAYER M2 ;
        RECT 15.31 30.52 16.51 30.8 ;
  LAYER M3 ;
        RECT 16.2 24.2 16.48 28.72 ;
  LAYER M3 ;
        RECT 15.77 24.62 16.05 29.14 ;
  LAYER M2 ;
        RECT 14.88 25.06 16.94 25.34 ;
  LAYER M1 ;
        RECT 16.215 16.295 16.465 19.825 ;
  LAYER M1 ;
        RECT 16.215 20.075 16.465 21.085 ;
  LAYER M1 ;
        RECT 16.215 22.175 16.465 23.185 ;
  LAYER M1 ;
        RECT 16.645 16.295 16.895 19.825 ;
  LAYER M1 ;
        RECT 15.785 16.295 16.035 19.825 ;
  LAYER M1 ;
        RECT 15.355 16.295 15.605 19.825 ;
  LAYER M1 ;
        RECT 15.355 20.075 15.605 21.085 ;
  LAYER M1 ;
        RECT 15.355 22.175 15.605 23.185 ;
  LAYER M1 ;
        RECT 14.925 16.295 15.175 19.825 ;
  LAYER M2 ;
        RECT 15.31 22.54 16.51 22.82 ;
  LAYER M2 ;
        RECT 16.17 16.24 17.37 16.52 ;
  LAYER M2 ;
        RECT 15.31 16.66 16.51 16.94 ;
  LAYER M2 ;
        RECT 16.17 20.44 17.37 20.72 ;
  LAYER M2 ;
        RECT 15.31 20.86 16.51 21.14 ;
  LAYER M2 ;
        RECT 14.88 17.08 16.94 17.36 ;
  LAYER M1 ;
        RECT 24.815 16.295 25.065 19.825 ;
  LAYER M1 ;
        RECT 24.815 20.075 25.065 21.085 ;
  LAYER M1 ;
        RECT 24.815 22.175 25.065 23.185 ;
  LAYER M1 ;
        RECT 18.795 16.295 19.045 19.825 ;
  LAYER M1 ;
        RECT 30.835 16.295 31.085 19.825 ;
  LAYER M2 ;
        RECT 24.34 16.24 25.54 16.52 ;
  LAYER M2 ;
        RECT 18.75 16.66 31.13 16.94 ;
  LAYER M2 ;
        RECT 24.34 22.54 25.54 22.82 ;
  LAYER M2 ;
        RECT 23.91 20.44 25.11 20.72 ;
  LAYER M3 ;
        RECT 25.23 16.22 25.51 22.84 ;
  LAYER M1 ;
        RECT 6.755 16.295 7.005 19.825 ;
  LAYER M1 ;
        RECT 6.755 20.075 7.005 21.085 ;
  LAYER M1 ;
        RECT 6.755 22.175 7.005 23.185 ;
  LAYER M1 ;
        RECT 12.775 16.295 13.025 19.825 ;
  LAYER M1 ;
        RECT 0.735 16.295 0.985 19.825 ;
  LAYER M2 ;
        RECT 6.28 16.24 7.48 16.52 ;
  LAYER M2 ;
        RECT 0.69 16.66 13.07 16.94 ;
  LAYER M2 ;
        RECT 6.28 22.54 7.48 22.82 ;
  LAYER M2 ;
        RECT 6.71 20.44 7.91 20.72 ;
  LAYER M3 ;
        RECT 6.31 16.22 6.59 22.84 ;
  LAYER M3 ;
        RECT 47.59 2.78 47.87 7.3 ;
  LAYER M2 ;
        RECT 46.7 10.78 47.9 11.06 ;
  LAYER M2 ;
        RECT 38.96 10.78 40.16 11.06 ;
  LAYER M3 ;
        RECT 47.59 7.14 47.87 10.92 ;
  LAYER M2 ;
        RECT 47.57 10.78 47.89 11.06 ;
  LAYER M2 ;
        RECT 39.99 10.78 46.87 11.06 ;
  LAYER M2 ;
        RECT 47.57 10.78 47.89 11.06 ;
  LAYER M3 ;
        RECT 47.59 10.76 47.87 11.08 ;
  LAYER M2 ;
        RECT 47.57 10.78 47.89 11.06 ;
  LAYER M3 ;
        RECT 47.59 10.76 47.87 11.08 ;
  LAYER M2 ;
        RECT 47.57 10.78 47.89 11.06 ;
  LAYER M3 ;
        RECT 47.59 10.76 47.87 11.08 ;
  LAYER M2 ;
        RECT 47.57 10.78 47.89 11.06 ;
  LAYER M3 ;
        RECT 47.59 10.76 47.87 11.08 ;
  LAYER M3 ;
        RECT 48.02 2.36 48.3 6.88 ;
  LAYER M2 ;
        RECT 47.56 10.36 48.76 10.64 ;
  LAYER M2 ;
        RECT 56.16 10.78 57.36 11.06 ;
  LAYER M3 ;
        RECT 48.02 6.72 48.3 10.5 ;
  LAYER M2 ;
        RECT 48 10.36 48.32 10.64 ;
  LAYER M2 ;
        RECT 48.43 10.36 48.75 10.64 ;
  LAYER M3 ;
        RECT 48.45 10.5 48.73 10.92 ;
  LAYER M2 ;
        RECT 48.59 10.78 56.33 11.06 ;
  LAYER M2 ;
        RECT 48 10.36 48.32 10.64 ;
  LAYER M3 ;
        RECT 48.02 10.34 48.3 10.66 ;
  LAYER M2 ;
        RECT 48 10.36 48.32 10.64 ;
  LAYER M3 ;
        RECT 48.02 10.34 48.3 10.66 ;
  LAYER M2 ;
        RECT 48.43 10.36 48.75 10.64 ;
  LAYER M3 ;
        RECT 48.45 10.34 48.73 10.66 ;
  LAYER M2 ;
        RECT 48.43 10.78 48.75 11.06 ;
  LAYER M3 ;
        RECT 48.45 10.76 48.73 11.08 ;
  LAYER M2 ;
        RECT 48 10.36 48.32 10.64 ;
  LAYER M3 ;
        RECT 48.02 10.34 48.3 10.66 ;
  LAYER M2 ;
        RECT 48.43 10.36 48.75 10.64 ;
  LAYER M3 ;
        RECT 48.45 10.34 48.73 10.66 ;
  LAYER M2 ;
        RECT 48.43 10.78 48.75 11.06 ;
  LAYER M3 ;
        RECT 48.45 10.76 48.73 11.08 ;
  LAYER M2 ;
        RECT 48 10.36 48.32 10.64 ;
  LAYER M3 ;
        RECT 48.02 10.34 48.3 10.66 ;
  LAYER M1 ;
        RECT 47.605 3.695 47.855 7.225 ;
  LAYER M1 ;
        RECT 47.605 2.435 47.855 3.445 ;
  LAYER M1 ;
        RECT 47.605 0.335 47.855 1.345 ;
  LAYER M1 ;
        RECT 47.175 3.695 47.425 7.225 ;
  LAYER M1 ;
        RECT 48.035 3.695 48.285 7.225 ;
  LAYER M1 ;
        RECT 48.465 3.695 48.715 7.225 ;
  LAYER M1 ;
        RECT 48.465 2.435 48.715 3.445 ;
  LAYER M1 ;
        RECT 48.465 0.335 48.715 1.345 ;
  LAYER M1 ;
        RECT 48.895 3.695 49.145 7.225 ;
  LAYER M2 ;
        RECT 46.7 7 47.9 7.28 ;
  LAYER M2 ;
        RECT 47.56 2.8 48.76 3.08 ;
  LAYER M2 ;
        RECT 47.56 6.58 48.76 6.86 ;
  LAYER M2 ;
        RECT 47.13 2.38 48.33 2.66 ;
  LAYER M2 ;
        RECT 47.56 0.7 48.76 0.98 ;
  LAYER M3 ;
        RECT 47.59 2.78 47.87 7.3 ;
  LAYER M3 ;
        RECT 48.02 2.36 48.3 6.88 ;
  LAYER M2 ;
        RECT 47.13 6.16 49.19 6.44 ;
  LAYER M1 ;
        RECT 47.605 11.675 47.855 15.205 ;
  LAYER M1 ;
        RECT 47.605 10.415 47.855 11.425 ;
  LAYER M1 ;
        RECT 47.605 8.315 47.855 9.325 ;
  LAYER M1 ;
        RECT 47.175 11.675 47.425 15.205 ;
  LAYER M1 ;
        RECT 48.035 11.675 48.285 15.205 ;
  LAYER M1 ;
        RECT 48.465 11.675 48.715 15.205 ;
  LAYER M1 ;
        RECT 48.465 10.415 48.715 11.425 ;
  LAYER M1 ;
        RECT 48.465 8.315 48.715 9.325 ;
  LAYER M1 ;
        RECT 48.895 11.675 49.145 15.205 ;
  LAYER M2 ;
        RECT 47.56 8.68 48.76 8.96 ;
  LAYER M2 ;
        RECT 46.7 14.98 47.9 15.26 ;
  LAYER M2 ;
        RECT 47.56 14.56 48.76 14.84 ;
  LAYER M2 ;
        RECT 46.7 10.78 47.9 11.06 ;
  LAYER M2 ;
        RECT 47.56 10.36 48.76 10.64 ;
  LAYER M2 ;
        RECT 47.13 14.14 49.19 14.42 ;
  LAYER M1 ;
        RECT 39.005 11.675 39.255 15.205 ;
  LAYER M1 ;
        RECT 39.005 10.415 39.255 11.425 ;
  LAYER M1 ;
        RECT 39.005 8.315 39.255 9.325 ;
  LAYER M1 ;
        RECT 45.025 11.675 45.275 15.205 ;
  LAYER M1 ;
        RECT 32.985 11.675 33.235 15.205 ;
  LAYER M2 ;
        RECT 38.53 14.98 39.73 15.26 ;
  LAYER M2 ;
        RECT 32.94 14.56 45.32 14.84 ;
  LAYER M2 ;
        RECT 38.53 8.68 39.73 8.96 ;
  LAYER M2 ;
        RECT 38.96 10.78 40.16 11.06 ;
  LAYER M3 ;
        RECT 38.56 8.66 38.84 15.28 ;
  LAYER M1 ;
        RECT 57.065 11.675 57.315 15.205 ;
  LAYER M1 ;
        RECT 57.065 10.415 57.315 11.425 ;
  LAYER M1 ;
        RECT 57.065 8.315 57.315 9.325 ;
  LAYER M1 ;
        RECT 51.045 11.675 51.295 15.205 ;
  LAYER M1 ;
        RECT 63.085 11.675 63.335 15.205 ;
  LAYER M2 ;
        RECT 56.59 14.98 57.79 15.26 ;
  LAYER M2 ;
        RECT 51 14.56 63.38 14.84 ;
  LAYER M2 ;
        RECT 56.59 8.68 57.79 8.96 ;
  LAYER M2 ;
        RECT 56.16 10.78 57.36 11.06 ;
  LAYER M3 ;
        RECT 57.48 8.66 57.76 15.28 ;
  LAYER M3 ;
        RECT 47.59 24.2 47.87 28.72 ;
  LAYER M2 ;
        RECT 46.7 20.44 47.9 20.72 ;
  LAYER M2 ;
        RECT 38.96 20.44 40.16 20.72 ;
  LAYER M3 ;
        RECT 47.59 20.58 47.87 24.36 ;
  LAYER M2 ;
        RECT 47.57 20.44 47.89 20.72 ;
  LAYER M2 ;
        RECT 39.99 20.44 46.87 20.72 ;
  LAYER M2 ;
        RECT 47.57 20.44 47.89 20.72 ;
  LAYER M3 ;
        RECT 47.59 20.42 47.87 20.74 ;
  LAYER M2 ;
        RECT 47.57 20.44 47.89 20.72 ;
  LAYER M3 ;
        RECT 47.59 20.42 47.87 20.74 ;
  LAYER M2 ;
        RECT 47.57 20.44 47.89 20.72 ;
  LAYER M3 ;
        RECT 47.59 20.42 47.87 20.74 ;
  LAYER M2 ;
        RECT 47.57 20.44 47.89 20.72 ;
  LAYER M3 ;
        RECT 47.59 20.42 47.87 20.74 ;
  LAYER M3 ;
        RECT 48.02 24.62 48.3 29.14 ;
  LAYER M2 ;
        RECT 47.56 20.86 48.76 21.14 ;
  LAYER M2 ;
        RECT 56.16 20.44 57.36 20.72 ;
  LAYER M3 ;
        RECT 48.02 21 48.3 24.78 ;
  LAYER M2 ;
        RECT 48 20.86 48.32 21.14 ;
  LAYER M2 ;
        RECT 48.43 20.86 48.75 21.14 ;
  LAYER M3 ;
        RECT 48.45 20.58 48.73 21 ;
  LAYER M2 ;
        RECT 48.59 20.44 56.33 20.72 ;
  LAYER M2 ;
        RECT 48 20.86 48.32 21.14 ;
  LAYER M3 ;
        RECT 48.02 20.84 48.3 21.16 ;
  LAYER M2 ;
        RECT 48 20.86 48.32 21.14 ;
  LAYER M3 ;
        RECT 48.02 20.84 48.3 21.16 ;
  LAYER M2 ;
        RECT 48.43 20.86 48.75 21.14 ;
  LAYER M3 ;
        RECT 48.45 20.84 48.73 21.16 ;
  LAYER M2 ;
        RECT 48.43 20.44 48.75 20.72 ;
  LAYER M3 ;
        RECT 48.45 20.42 48.73 20.74 ;
  LAYER M2 ;
        RECT 48 20.86 48.32 21.14 ;
  LAYER M3 ;
        RECT 48.02 20.84 48.3 21.16 ;
  LAYER M2 ;
        RECT 48.43 20.86 48.75 21.14 ;
  LAYER M3 ;
        RECT 48.45 20.84 48.73 21.16 ;
  LAYER M2 ;
        RECT 48.43 20.44 48.75 20.72 ;
  LAYER M3 ;
        RECT 48.45 20.42 48.73 20.74 ;
  LAYER M2 ;
        RECT 48 20.86 48.32 21.14 ;
  LAYER M3 ;
        RECT 48.02 20.84 48.3 21.16 ;
  LAYER M1 ;
        RECT 47.605 24.275 47.855 27.805 ;
  LAYER M1 ;
        RECT 47.605 28.055 47.855 29.065 ;
  LAYER M1 ;
        RECT 47.605 30.155 47.855 31.165 ;
  LAYER M1 ;
        RECT 47.175 24.275 47.425 27.805 ;
  LAYER M1 ;
        RECT 48.035 24.275 48.285 27.805 ;
  LAYER M1 ;
        RECT 48.465 24.275 48.715 27.805 ;
  LAYER M1 ;
        RECT 48.465 28.055 48.715 29.065 ;
  LAYER M1 ;
        RECT 48.465 30.155 48.715 31.165 ;
  LAYER M1 ;
        RECT 48.895 24.275 49.145 27.805 ;
  LAYER M2 ;
        RECT 46.7 24.22 47.9 24.5 ;
  LAYER M2 ;
        RECT 47.56 28.42 48.76 28.7 ;
  LAYER M2 ;
        RECT 47.56 24.64 48.76 24.92 ;
  LAYER M2 ;
        RECT 47.13 28.84 48.33 29.12 ;
  LAYER M2 ;
        RECT 47.56 30.52 48.76 30.8 ;
  LAYER M3 ;
        RECT 47.59 24.2 47.87 28.72 ;
  LAYER M3 ;
        RECT 48.02 24.62 48.3 29.14 ;
  LAYER M2 ;
        RECT 47.13 25.06 49.19 25.34 ;
  LAYER M1 ;
        RECT 47.605 16.295 47.855 19.825 ;
  LAYER M1 ;
        RECT 47.605 20.075 47.855 21.085 ;
  LAYER M1 ;
        RECT 47.605 22.175 47.855 23.185 ;
  LAYER M1 ;
        RECT 47.175 16.295 47.425 19.825 ;
  LAYER M1 ;
        RECT 48.035 16.295 48.285 19.825 ;
  LAYER M1 ;
        RECT 48.465 16.295 48.715 19.825 ;
  LAYER M1 ;
        RECT 48.465 20.075 48.715 21.085 ;
  LAYER M1 ;
        RECT 48.465 22.175 48.715 23.185 ;
  LAYER M1 ;
        RECT 48.895 16.295 49.145 19.825 ;
  LAYER M2 ;
        RECT 47.56 22.54 48.76 22.82 ;
  LAYER M2 ;
        RECT 46.7 16.24 47.9 16.52 ;
  LAYER M2 ;
        RECT 47.56 16.66 48.76 16.94 ;
  LAYER M2 ;
        RECT 46.7 20.44 47.9 20.72 ;
  LAYER M2 ;
        RECT 47.56 20.86 48.76 21.14 ;
  LAYER M2 ;
        RECT 47.13 17.08 49.19 17.36 ;
  LAYER M1 ;
        RECT 39.005 16.295 39.255 19.825 ;
  LAYER M1 ;
        RECT 39.005 20.075 39.255 21.085 ;
  LAYER M1 ;
        RECT 39.005 22.175 39.255 23.185 ;
  LAYER M1 ;
        RECT 45.025 16.295 45.275 19.825 ;
  LAYER M1 ;
        RECT 32.985 16.295 33.235 19.825 ;
  LAYER M2 ;
        RECT 38.53 16.24 39.73 16.52 ;
  LAYER M2 ;
        RECT 32.94 16.66 45.32 16.94 ;
  LAYER M2 ;
        RECT 38.53 22.54 39.73 22.82 ;
  LAYER M2 ;
        RECT 38.96 20.44 40.16 20.72 ;
  LAYER M3 ;
        RECT 38.56 16.22 38.84 22.84 ;
  LAYER M1 ;
        RECT 57.065 16.295 57.315 19.825 ;
  LAYER M1 ;
        RECT 57.065 20.075 57.315 21.085 ;
  LAYER M1 ;
        RECT 57.065 22.175 57.315 23.185 ;
  LAYER M1 ;
        RECT 51.045 16.295 51.295 19.825 ;
  LAYER M1 ;
        RECT 63.085 16.295 63.335 19.825 ;
  LAYER M2 ;
        RECT 56.59 16.24 57.79 16.52 ;
  LAYER M2 ;
        RECT 51 16.66 63.38 16.94 ;
  LAYER M2 ;
        RECT 56.59 22.54 57.79 22.82 ;
  LAYER M2 ;
        RECT 56.16 20.44 57.36 20.72 ;
  LAYER M3 ;
        RECT 57.48 16.22 57.76 22.84 ;
  END 
END DCDC_CONV2TO1_1
