MACRO CCP_NMOS_B_26073270_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CCP_NMOS_B_26073270_X1_Y1 0 0 ;
  SIZE 5160 BY 9240 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1980 7420 3180 7700 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2010 1100 2290 5620 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2440 1520 2720 6040 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1550 1960 3610 2240 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 2025 1175 2275 4705 ;
    LAYER M1 ;
      RECT 2025 4955 2275 5965 ;
    LAYER M1 ;
      RECT 2025 7055 2275 8065 ;
    LAYER M1 ;
      RECT 1595 1175 1845 4705 ;
    LAYER M1 ;
      RECT 2455 1175 2705 4705 ;
    LAYER M1 ;
      RECT 2885 1175 3135 4705 ;
    LAYER M1 ;
      RECT 2885 4955 3135 5965 ;
    LAYER M1 ;
      RECT 2885 7055 3135 8065 ;
    LAYER M1 ;
      RECT 3315 1175 3565 4705 ;
    LAYER M2 ;
      RECT 1120 1120 2320 1400 ;
    LAYER M2 ;
      RECT 1980 5320 3180 5600 ;
    LAYER M2 ;
      RECT 1980 1540 3180 1820 ;
    LAYER M2 ;
      RECT 1550 5740 2750 6020 ;
    LAYER V1 ;
      RECT 2065 1175 2235 1345 ;
    LAYER V1 ;
      RECT 2065 5795 2235 5965 ;
    LAYER V1 ;
      RECT 2065 7475 2235 7645 ;
    LAYER V1 ;
      RECT 2925 1595 3095 1765 ;
    LAYER V1 ;
      RECT 2925 5375 3095 5545 ;
    LAYER V1 ;
      RECT 2925 7475 3095 7645 ;
    LAYER V1 ;
      RECT 1635 2015 1805 2185 ;
    LAYER V1 ;
      RECT 2495 2015 2665 2185 ;
    LAYER V1 ;
      RECT 3355 2015 3525 2185 ;
    LAYER V2 ;
      RECT 2075 1185 2225 1335 ;
    LAYER V2 ;
      RECT 2075 5385 2225 5535 ;
    LAYER V2 ;
      RECT 2505 1605 2655 1755 ;
    LAYER V2 ;
      RECT 2505 5805 2655 5955 ;
    LAYER V0 ;
      RECT 2065 3545 2235 3715 ;
    LAYER V0 ;
      RECT 2065 5375 2235 5545 ;
    LAYER V0 ;
      RECT 2065 7475 2235 7645 ;
    LAYER V0 ;
      RECT 1635 3545 1805 3715 ;
    LAYER V0 ;
      RECT 2495 3545 2665 3715 ;
    LAYER V0 ;
      RECT 2495 3545 2665 3715 ;
    LAYER V0 ;
      RECT 2925 3545 3095 3715 ;
    LAYER V0 ;
      RECT 2925 5375 3095 5545 ;
    LAYER V0 ;
      RECT 2925 7475 3095 7645 ;
    LAYER V0 ;
      RECT 3355 3545 3525 3715 ;
  END
END CCP_NMOS_B_26073270_X1_Y1
