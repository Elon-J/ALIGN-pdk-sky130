MACRO DCDC_CONV2TO1_1
  ORIGIN 0 0 ;
  FOREIGN DCDC_CONV2TO1_1 0 0 ;
  SIZE 61.92 BY 30.24 ;
  PIN CLK0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 6.31 15.38 6.59 22 ;
      LAYER M3 ;
        RECT 55.33 15.38 55.61 22 ;
      LAYER M3 ;
        RECT 6.31 16.195 6.59 16.565 ;
      LAYER M4 ;
        RECT 6.45 15.98 55.47 16.78 ;
      LAYER M3 ;
        RECT 55.33 16.195 55.61 16.565 ;
    END
  END CLK0
  PIN CLK0B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 24.37 8.24 24.65 14.86 ;
      LAYER M3 ;
        RECT 37.27 8.24 37.55 14.86 ;
      LAYER M3 ;
        RECT 24.37 7.98 24.65 8.4 ;
      LAYER M2 ;
        RECT 24.51 7.84 37.41 8.12 ;
      LAYER M3 ;
        RECT 37.27 7.98 37.55 8.4 ;
    END
  END CLK0B
  PIN CLK1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 24.37 15.38 24.65 22 ;
      LAYER M3 ;
        RECT 37.27 15.38 37.55 22 ;
      LAYER M3 ;
        RECT 24.37 21.84 24.65 22.68 ;
      LAYER M4 ;
        RECT 24.51 22.28 25.16 23.08 ;
      LAYER M5 ;
        RECT 24.57 22.68 25.75 25.2 ;
      LAYER M4 ;
        RECT 25.16 24.8 37 25.6 ;
      LAYER M5 ;
        RECT 36.41 23.94 37.59 25.2 ;
      LAYER M4 ;
        RECT 37 23.54 37.41 24.34 ;
      LAYER M3 ;
        RECT 37.27 21.84 37.55 23.94 ;
    END
  END CLK1
  PIN CLK1B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 6.31 8.24 6.59 14.86 ;
      LAYER M3 ;
        RECT 55.33 8.24 55.61 14.86 ;
      LAYER M3 ;
        RECT 6.31 11.155 6.59 11.525 ;
      LAYER M4 ;
        RECT 6.45 10.94 55.47 11.74 ;
      LAYER M3 ;
        RECT 55.33 11.155 55.61 11.525 ;
    END
  END CLK1B
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.88 29.26 16.08 29.54 ;
      LAYER M2 ;
        RECT 14.88 21.7 16.08 21.98 ;
      LAYER M2 ;
        RECT 14.89 29.26 15.21 29.54 ;
      LAYER M3 ;
        RECT 14.91 21.84 15.19 29.4 ;
      LAYER M2 ;
        RECT 14.89 21.7 15.21 21.98 ;
      LAYER M2 ;
        RECT 45.84 29.26 47.04 29.54 ;
      LAYER M2 ;
        RECT 45.84 21.7 47.04 21.98 ;
      LAYER M2 ;
        RECT 46.71 29.26 47.03 29.54 ;
      LAYER M3 ;
        RECT 46.73 21.84 47.01 29.4 ;
      LAYER M2 ;
        RECT 46.71 21.7 47.03 21.98 ;
      LAYER M2 ;
        RECT 15.91 21.7 16.34 21.98 ;
      LAYER M3 ;
        RECT 16.2 21.42 16.48 21.84 ;
      LAYER M4 ;
        RECT 16.34 21.02 43 21.82 ;
      LAYER M3 ;
        RECT 42.86 21.42 43.14 21.84 ;
      LAYER M2 ;
        RECT 43 21.7 46.01 21.98 ;
    END
  END VGND
  PIN VHIGH
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.45 6.16 16.51 6.44 ;
      LAYER M2 ;
        RECT 14.45 13.72 16.51 14 ;
      LAYER M2 ;
        RECT 14.46 6.16 14.78 6.44 ;
      LAYER M3 ;
        RECT 14.48 6.3 14.76 13.86 ;
      LAYER M2 ;
        RECT 14.46 13.72 14.78 14 ;
    END
  END VHIGH
  PIN VMID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.45 23.8 16.51 24.08 ;
      LAYER M2 ;
        RECT 14.45 16.24 16.51 16.52 ;
      LAYER M2 ;
        RECT 14.46 23.8 14.78 24.08 ;
      LAYER M3 ;
        RECT 14.48 16.38 14.76 23.94 ;
      LAYER M2 ;
        RECT 14.46 16.24 14.78 16.52 ;
      LAYER M2 ;
        RECT 45.41 6.16 47.47 6.44 ;
      LAYER M2 ;
        RECT 45.41 13.72 47.47 14 ;
      LAYER M2 ;
        RECT 45.42 6.16 45.74 6.44 ;
      LAYER M3 ;
        RECT 45.44 6.3 45.72 13.86 ;
      LAYER M2 ;
        RECT 45.42 13.72 45.74 14 ;
      LAYER M2 ;
        RECT 16.34 16.24 17.2 16.52 ;
      LAYER M1 ;
        RECT 17.075 13.86 17.325 16.38 ;
      LAYER M2 ;
        RECT 17.2 13.72 45.58 14 ;
    END
  END VMID
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.88 0.7 16.08 0.98 ;
      LAYER M2 ;
        RECT 14.88 8.26 16.08 8.54 ;
      LAYER M2 ;
        RECT 14.89 0.7 15.21 0.98 ;
      LAYER M3 ;
        RECT 14.91 0.84 15.19 8.4 ;
      LAYER M2 ;
        RECT 14.89 8.26 15.21 8.54 ;
      LAYER M2 ;
        RECT 45.84 0.7 47.04 0.98 ;
      LAYER M2 ;
        RECT 45.84 8.26 47.04 8.54 ;
      LAYER M2 ;
        RECT 46.71 0.7 47.03 0.98 ;
      LAYER M3 ;
        RECT 46.73 0.84 47.01 8.4 ;
      LAYER M2 ;
        RECT 46.71 8.26 47.03 8.54 ;
      LAYER M2 ;
        RECT 15.75 0.7 16.07 0.98 ;
      LAYER M3 ;
        RECT 15.77 0.84 16.05 1.26 ;
      LAYER M4 ;
        RECT 15.91 0.86 43 1.66 ;
      LAYER M3 ;
        RECT 42.86 0.84 43.14 1.26 ;
      LAYER M2 ;
        RECT 43 0.7 46.01 0.98 ;
    END
  END VPWR
  PIN Y0_TOP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.74 14.56 16.94 14.84 ;
      LAYER M2 ;
        RECT 15.74 15.4 16.94 15.68 ;
      LAYER M2 ;
        RECT 16.18 14.56 16.5 14.84 ;
      LAYER M3 ;
        RECT 16.2 14.7 16.48 15.54 ;
      LAYER M2 ;
        RECT 16.18 15.4 16.5 15.68 ;
    END
  END Y0_TOP
  PIN Y1_TOP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.88 14.14 16.08 14.42 ;
      LAYER M2 ;
        RECT 14.88 15.82 16.08 16.1 ;
      LAYER M2 ;
        RECT 15.32 14.14 15.64 14.42 ;
      LAYER M3 ;
        RECT 15.34 14.28 15.62 15.96 ;
      LAYER M2 ;
        RECT 15.32 15.82 15.64 16.1 ;
    END
  END Y1_TOP
  PIN VLOW
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 45.41 23.8 47.47 24.08 ;
      LAYER M2 ;
        RECT 45.41 16.24 47.47 16.52 ;
      LAYER M2 ;
        RECT 45.42 23.8 45.74 24.08 ;
      LAYER M3 ;
        RECT 45.44 16.38 45.72 23.94 ;
      LAYER M2 ;
        RECT 45.42 16.24 45.74 16.52 ;
    END
  END VLOW
  PIN Y0_BOT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 44.98 14.56 46.18 14.84 ;
      LAYER M2 ;
        RECT 44.98 15.4 46.18 15.68 ;
      LAYER M2 ;
        RECT 45.42 14.56 45.74 14.84 ;
      LAYER M3 ;
        RECT 45.44 14.7 45.72 15.54 ;
      LAYER M2 ;
        RECT 45.42 15.4 45.74 15.68 ;
    END
  END Y0_BOT
  PIN Y1_BOT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 45.84 14.14 47.04 14.42 ;
      LAYER M2 ;
        RECT 45.84 15.82 47.04 16.1 ;
      LAYER M2 ;
        RECT 46.28 14.14 46.6 14.42 ;
      LAYER M3 ;
        RECT 46.3 14.28 46.58 15.96 ;
      LAYER M2 ;
        RECT 46.28 15.82 46.6 16.1 ;
    END
  END Y1_BOT
  OBS 
  LAYER M3 ;
        RECT 15.77 2.78 16.05 7.3 ;
  LAYER M2 ;
        RECT 15.74 10.36 16.94 10.64 ;
  LAYER M2 ;
        RECT 23.05 10.36 24.25 10.64 ;
  LAYER M3 ;
        RECT 15.77 7.14 16.05 10.5 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M2 ;
        RECT 16.77 10.36 23.22 10.64 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M3 ;
        RECT 15.34 2.36 15.62 6.88 ;
  LAYER M2 ;
        RECT 14.88 9.94 16.08 10.22 ;
  LAYER M2 ;
        RECT 6.71 10.36 7.91 10.64 ;
  LAYER M3 ;
        RECT 15.34 6.72 15.62 10.08 ;
  LAYER M2 ;
        RECT 15.32 9.94 15.64 10.22 ;
  LAYER M2 ;
        RECT 14.89 9.94 15.21 10.22 ;
  LAYER M3 ;
        RECT 14.91 10.08 15.19 10.5 ;
  LAYER M2 ;
        RECT 7.74 10.36 15.05 10.64 ;
  LAYER M2 ;
        RECT 15.32 9.94 15.64 10.22 ;
  LAYER M3 ;
        RECT 15.34 9.92 15.62 10.24 ;
  LAYER M2 ;
        RECT 15.32 9.94 15.64 10.22 ;
  LAYER M3 ;
        RECT 15.34 9.92 15.62 10.24 ;
  LAYER M2 ;
        RECT 14.89 9.94 15.21 10.22 ;
  LAYER M3 ;
        RECT 14.91 9.92 15.19 10.24 ;
  LAYER M2 ;
        RECT 14.89 10.36 15.21 10.64 ;
  LAYER M3 ;
        RECT 14.91 10.34 15.19 10.66 ;
  LAYER M2 ;
        RECT 15.32 9.94 15.64 10.22 ;
  LAYER M3 ;
        RECT 15.34 9.92 15.62 10.24 ;
  LAYER M2 ;
        RECT 14.89 9.94 15.21 10.22 ;
  LAYER M3 ;
        RECT 14.91 9.92 15.19 10.24 ;
  LAYER M2 ;
        RECT 14.89 10.36 15.21 10.64 ;
  LAYER M3 ;
        RECT 14.91 10.34 15.19 10.66 ;
  LAYER M2 ;
        RECT 15.32 9.94 15.64 10.22 ;
  LAYER M3 ;
        RECT 15.34 9.92 15.62 10.24 ;
  LAYER M1 ;
        RECT 15.785 3.695 16.035 7.225 ;
  LAYER M1 ;
        RECT 15.785 2.435 16.035 3.445 ;
  LAYER M1 ;
        RECT 15.785 0.335 16.035 1.345 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M1 ;
        RECT 14.925 2.435 15.175 3.445 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 1.345 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M2 ;
        RECT 15.74 7 16.94 7.28 ;
  LAYER M2 ;
        RECT 14.88 2.8 16.08 3.08 ;
  LAYER M2 ;
        RECT 14.88 6.58 16.08 6.86 ;
  LAYER M2 ;
        RECT 15.31 2.38 16.51 2.66 ;
  LAYER M2 ;
        RECT 14.88 0.7 16.08 0.98 ;
  LAYER M3 ;
        RECT 15.77 2.78 16.05 7.3 ;
  LAYER M3 ;
        RECT 15.34 2.36 15.62 6.88 ;
  LAYER M2 ;
        RECT 14.45 6.16 16.51 6.44 ;
  LAYER M1 ;
        RECT 15.785 11.255 16.035 14.785 ;
  LAYER M1 ;
        RECT 15.785 9.995 16.035 11.005 ;
  LAYER M1 ;
        RECT 15.785 7.895 16.035 8.905 ;
  LAYER M1 ;
        RECT 16.215 11.255 16.465 14.785 ;
  LAYER M1 ;
        RECT 15.355 11.255 15.605 14.785 ;
  LAYER M1 ;
        RECT 14.925 11.255 15.175 14.785 ;
  LAYER M1 ;
        RECT 14.925 9.995 15.175 11.005 ;
  LAYER M1 ;
        RECT 14.925 7.895 15.175 8.905 ;
  LAYER M1 ;
        RECT 14.495 11.255 14.745 14.785 ;
  LAYER M2 ;
        RECT 14.88 8.26 16.08 8.54 ;
  LAYER M2 ;
        RECT 15.74 14.56 16.94 14.84 ;
  LAYER M2 ;
        RECT 14.88 14.14 16.08 14.42 ;
  LAYER M2 ;
        RECT 15.74 10.36 16.94 10.64 ;
  LAYER M2 ;
        RECT 14.88 9.94 16.08 10.22 ;
  LAYER M2 ;
        RECT 14.45 13.72 16.51 14 ;
  LAYER M1 ;
        RECT 23.955 11.255 24.205 14.785 ;
  LAYER M1 ;
        RECT 23.955 9.995 24.205 11.005 ;
  LAYER M1 ;
        RECT 23.955 7.895 24.205 8.905 ;
  LAYER M1 ;
        RECT 17.935 11.255 18.185 14.785 ;
  LAYER M1 ;
        RECT 29.975 11.255 30.225 14.785 ;
  LAYER M2 ;
        RECT 17.89 14.56 30.27 14.84 ;
  LAYER M2 ;
        RECT 23.48 8.26 24.68 8.54 ;
  LAYER M2 ;
        RECT 23.48 14.14 24.68 14.42 ;
  LAYER M2 ;
        RECT 23.05 10.36 24.25 10.64 ;
  LAYER M3 ;
        RECT 24.37 8.24 24.65 14.86 ;
  LAYER M1 ;
        RECT 6.755 11.255 7.005 14.785 ;
  LAYER M1 ;
        RECT 6.755 9.995 7.005 11.005 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 8.905 ;
  LAYER M1 ;
        RECT 12.775 11.255 13.025 14.785 ;
  LAYER M1 ;
        RECT 0.735 11.255 0.985 14.785 ;
  LAYER M2 ;
        RECT 0.69 14.56 13.07 14.84 ;
  LAYER M2 ;
        RECT 6.28 8.26 7.48 8.54 ;
  LAYER M2 ;
        RECT 6.28 14.14 7.48 14.42 ;
  LAYER M2 ;
        RECT 6.71 10.36 7.91 10.64 ;
  LAYER M3 ;
        RECT 6.31 8.24 6.59 14.86 ;
  LAYER M3 ;
        RECT 15.77 22.94 16.05 27.46 ;
  LAYER M2 ;
        RECT 15.74 19.6 16.94 19.88 ;
  LAYER M2 ;
        RECT 23.05 19.6 24.25 19.88 ;
  LAYER M3 ;
        RECT 15.77 19.74 16.05 23.1 ;
  LAYER M2 ;
        RECT 15.75 19.6 16.07 19.88 ;
  LAYER M2 ;
        RECT 16.77 19.6 23.22 19.88 ;
  LAYER M2 ;
        RECT 15.75 19.6 16.07 19.88 ;
  LAYER M3 ;
        RECT 15.77 19.58 16.05 19.9 ;
  LAYER M2 ;
        RECT 15.75 19.6 16.07 19.88 ;
  LAYER M3 ;
        RECT 15.77 19.58 16.05 19.9 ;
  LAYER M2 ;
        RECT 15.75 19.6 16.07 19.88 ;
  LAYER M3 ;
        RECT 15.77 19.58 16.05 19.9 ;
  LAYER M2 ;
        RECT 15.75 19.6 16.07 19.88 ;
  LAYER M3 ;
        RECT 15.77 19.58 16.05 19.9 ;
  LAYER M3 ;
        RECT 15.34 23.36 15.62 27.88 ;
  LAYER M2 ;
        RECT 14.88 20.02 16.08 20.3 ;
  LAYER M2 ;
        RECT 6.71 19.6 7.91 19.88 ;
  LAYER M3 ;
        RECT 15.34 20.16 15.62 23.52 ;
  LAYER M2 ;
        RECT 15.32 20.02 15.64 20.3 ;
  LAYER M2 ;
        RECT 14.89 20.02 15.21 20.3 ;
  LAYER M3 ;
        RECT 14.91 19.74 15.19 20.16 ;
  LAYER M2 ;
        RECT 7.74 19.6 15.05 19.88 ;
  LAYER M2 ;
        RECT 15.32 20.02 15.64 20.3 ;
  LAYER M3 ;
        RECT 15.34 20 15.62 20.32 ;
  LAYER M2 ;
        RECT 15.32 20.02 15.64 20.3 ;
  LAYER M3 ;
        RECT 15.34 20 15.62 20.32 ;
  LAYER M2 ;
        RECT 14.89 19.6 15.21 19.88 ;
  LAYER M3 ;
        RECT 14.91 19.58 15.19 19.9 ;
  LAYER M2 ;
        RECT 14.89 20.02 15.21 20.3 ;
  LAYER M3 ;
        RECT 14.91 20 15.19 20.32 ;
  LAYER M2 ;
        RECT 15.32 20.02 15.64 20.3 ;
  LAYER M3 ;
        RECT 15.34 20 15.62 20.32 ;
  LAYER M2 ;
        RECT 14.89 19.6 15.21 19.88 ;
  LAYER M3 ;
        RECT 14.91 19.58 15.19 19.9 ;
  LAYER M2 ;
        RECT 14.89 20.02 15.21 20.3 ;
  LAYER M3 ;
        RECT 14.91 20 15.19 20.32 ;
  LAYER M2 ;
        RECT 15.32 20.02 15.64 20.3 ;
  LAYER M3 ;
        RECT 15.34 20 15.62 20.32 ;
  LAYER M1 ;
        RECT 15.785 23.015 16.035 26.545 ;
  LAYER M1 ;
        RECT 15.785 26.795 16.035 27.805 ;
  LAYER M1 ;
        RECT 15.785 28.895 16.035 29.905 ;
  LAYER M1 ;
        RECT 16.215 23.015 16.465 26.545 ;
  LAYER M1 ;
        RECT 15.355 23.015 15.605 26.545 ;
  LAYER M1 ;
        RECT 14.925 23.015 15.175 26.545 ;
  LAYER M1 ;
        RECT 14.925 26.795 15.175 27.805 ;
  LAYER M1 ;
        RECT 14.925 28.895 15.175 29.905 ;
  LAYER M1 ;
        RECT 14.495 23.015 14.745 26.545 ;
  LAYER M2 ;
        RECT 15.74 22.96 16.94 23.24 ;
  LAYER M2 ;
        RECT 14.88 27.16 16.08 27.44 ;
  LAYER M2 ;
        RECT 14.88 23.38 16.08 23.66 ;
  LAYER M2 ;
        RECT 15.31 27.58 16.51 27.86 ;
  LAYER M2 ;
        RECT 14.88 29.26 16.08 29.54 ;
  LAYER M3 ;
        RECT 15.77 22.94 16.05 27.46 ;
  LAYER M3 ;
        RECT 15.34 23.36 15.62 27.88 ;
  LAYER M2 ;
        RECT 14.45 23.8 16.51 24.08 ;
  LAYER M1 ;
        RECT 15.785 15.455 16.035 18.985 ;
  LAYER M1 ;
        RECT 15.785 19.235 16.035 20.245 ;
  LAYER M1 ;
        RECT 15.785 21.335 16.035 22.345 ;
  LAYER M1 ;
        RECT 16.215 15.455 16.465 18.985 ;
  LAYER M1 ;
        RECT 15.355 15.455 15.605 18.985 ;
  LAYER M1 ;
        RECT 14.925 15.455 15.175 18.985 ;
  LAYER M1 ;
        RECT 14.925 19.235 15.175 20.245 ;
  LAYER M1 ;
        RECT 14.925 21.335 15.175 22.345 ;
  LAYER M1 ;
        RECT 14.495 15.455 14.745 18.985 ;
  LAYER M2 ;
        RECT 14.88 21.7 16.08 21.98 ;
  LAYER M2 ;
        RECT 15.74 15.4 16.94 15.68 ;
  LAYER M2 ;
        RECT 14.88 15.82 16.08 16.1 ;
  LAYER M2 ;
        RECT 15.74 19.6 16.94 19.88 ;
  LAYER M2 ;
        RECT 14.88 20.02 16.08 20.3 ;
  LAYER M2 ;
        RECT 14.45 16.24 16.51 16.52 ;
  LAYER M1 ;
        RECT 23.955 15.455 24.205 18.985 ;
  LAYER M1 ;
        RECT 23.955 19.235 24.205 20.245 ;
  LAYER M1 ;
        RECT 23.955 21.335 24.205 22.345 ;
  LAYER M1 ;
        RECT 17.935 15.455 18.185 18.985 ;
  LAYER M1 ;
        RECT 29.975 15.455 30.225 18.985 ;
  LAYER M2 ;
        RECT 17.89 15.4 30.27 15.68 ;
  LAYER M2 ;
        RECT 23.48 21.7 24.68 21.98 ;
  LAYER M2 ;
        RECT 23.48 15.82 24.68 16.1 ;
  LAYER M2 ;
        RECT 23.05 19.6 24.25 19.88 ;
  LAYER M3 ;
        RECT 24.37 15.38 24.65 22 ;
  LAYER M1 ;
        RECT 6.755 15.455 7.005 18.985 ;
  LAYER M1 ;
        RECT 6.755 19.235 7.005 20.245 ;
  LAYER M1 ;
        RECT 6.755 21.335 7.005 22.345 ;
  LAYER M1 ;
        RECT 12.775 15.455 13.025 18.985 ;
  LAYER M1 ;
        RECT 0.735 15.455 0.985 18.985 ;
  LAYER M2 ;
        RECT 0.69 15.4 13.07 15.68 ;
  LAYER M2 ;
        RECT 6.28 21.7 7.48 21.98 ;
  LAYER M2 ;
        RECT 6.28 15.82 7.48 16.1 ;
  LAYER M2 ;
        RECT 6.71 19.6 7.91 19.88 ;
  LAYER M3 ;
        RECT 6.31 15.38 6.59 22 ;
  LAYER M3 ;
        RECT 45.87 2.78 46.15 7.3 ;
  LAYER M2 ;
        RECT 44.98 10.36 46.18 10.64 ;
  LAYER M2 ;
        RECT 37.67 10.36 38.87 10.64 ;
  LAYER M3 ;
        RECT 45.87 7.14 46.15 10.5 ;
  LAYER M2 ;
        RECT 45.85 10.36 46.17 10.64 ;
  LAYER M2 ;
        RECT 38.7 10.36 45.15 10.64 ;
  LAYER M2 ;
        RECT 45.85 10.36 46.17 10.64 ;
  LAYER M3 ;
        RECT 45.87 10.34 46.15 10.66 ;
  LAYER M2 ;
        RECT 45.85 10.36 46.17 10.64 ;
  LAYER M3 ;
        RECT 45.87 10.34 46.15 10.66 ;
  LAYER M2 ;
        RECT 45.85 10.36 46.17 10.64 ;
  LAYER M3 ;
        RECT 45.87 10.34 46.15 10.66 ;
  LAYER M2 ;
        RECT 45.85 10.36 46.17 10.64 ;
  LAYER M3 ;
        RECT 45.87 10.34 46.15 10.66 ;
  LAYER M3 ;
        RECT 46.3 2.36 46.58 6.88 ;
  LAYER M2 ;
        RECT 45.84 9.94 47.04 10.22 ;
  LAYER M2 ;
        RECT 54.01 10.36 55.21 10.64 ;
  LAYER M3 ;
        RECT 46.3 6.72 46.58 10.08 ;
  LAYER M2 ;
        RECT 46.28 9.94 46.6 10.22 ;
  LAYER M2 ;
        RECT 46.71 9.94 47.03 10.22 ;
  LAYER M3 ;
        RECT 46.73 10.08 47.01 10.5 ;
  LAYER M2 ;
        RECT 46.87 10.36 54.18 10.64 ;
  LAYER M2 ;
        RECT 46.28 9.94 46.6 10.22 ;
  LAYER M3 ;
        RECT 46.3 9.92 46.58 10.24 ;
  LAYER M2 ;
        RECT 46.28 9.94 46.6 10.22 ;
  LAYER M3 ;
        RECT 46.3 9.92 46.58 10.24 ;
  LAYER M2 ;
        RECT 46.28 9.94 46.6 10.22 ;
  LAYER M3 ;
        RECT 46.3 9.92 46.58 10.24 ;
  LAYER M2 ;
        RECT 46.71 9.94 47.03 10.22 ;
  LAYER M3 ;
        RECT 46.73 9.92 47.01 10.24 ;
  LAYER M2 ;
        RECT 46.71 10.36 47.03 10.64 ;
  LAYER M3 ;
        RECT 46.73 10.34 47.01 10.66 ;
  LAYER M2 ;
        RECT 46.28 9.94 46.6 10.22 ;
  LAYER M3 ;
        RECT 46.3 9.92 46.58 10.24 ;
  LAYER M2 ;
        RECT 46.71 9.94 47.03 10.22 ;
  LAYER M3 ;
        RECT 46.73 9.92 47.01 10.24 ;
  LAYER M2 ;
        RECT 46.71 10.36 47.03 10.64 ;
  LAYER M3 ;
        RECT 46.73 10.34 47.01 10.66 ;
  LAYER M1 ;
        RECT 45.885 3.695 46.135 7.225 ;
  LAYER M1 ;
        RECT 45.885 2.435 46.135 3.445 ;
  LAYER M1 ;
        RECT 45.885 0.335 46.135 1.345 ;
  LAYER M1 ;
        RECT 45.455 3.695 45.705 7.225 ;
  LAYER M1 ;
        RECT 46.315 3.695 46.565 7.225 ;
  LAYER M1 ;
        RECT 46.745 3.695 46.995 7.225 ;
  LAYER M1 ;
        RECT 46.745 2.435 46.995 3.445 ;
  LAYER M1 ;
        RECT 46.745 0.335 46.995 1.345 ;
  LAYER M1 ;
        RECT 47.175 3.695 47.425 7.225 ;
  LAYER M2 ;
        RECT 44.98 7 46.18 7.28 ;
  LAYER M2 ;
        RECT 45.84 2.8 47.04 3.08 ;
  LAYER M2 ;
        RECT 45.84 6.58 47.04 6.86 ;
  LAYER M2 ;
        RECT 45.41 2.38 46.61 2.66 ;
  LAYER M2 ;
        RECT 45.84 0.7 47.04 0.98 ;
  LAYER M3 ;
        RECT 45.87 2.78 46.15 7.3 ;
  LAYER M3 ;
        RECT 46.3 2.36 46.58 6.88 ;
  LAYER M2 ;
        RECT 45.41 6.16 47.47 6.44 ;
  LAYER M1 ;
        RECT 45.885 11.255 46.135 14.785 ;
  LAYER M1 ;
        RECT 45.885 9.995 46.135 11.005 ;
  LAYER M1 ;
        RECT 45.885 7.895 46.135 8.905 ;
  LAYER M1 ;
        RECT 45.455 11.255 45.705 14.785 ;
  LAYER M1 ;
        RECT 46.315 11.255 46.565 14.785 ;
  LAYER M1 ;
        RECT 46.745 11.255 46.995 14.785 ;
  LAYER M1 ;
        RECT 46.745 9.995 46.995 11.005 ;
  LAYER M1 ;
        RECT 46.745 7.895 46.995 8.905 ;
  LAYER M1 ;
        RECT 47.175 11.255 47.425 14.785 ;
  LAYER M2 ;
        RECT 45.84 8.26 47.04 8.54 ;
  LAYER M2 ;
        RECT 44.98 14.56 46.18 14.84 ;
  LAYER M2 ;
        RECT 45.84 14.14 47.04 14.42 ;
  LAYER M2 ;
        RECT 44.98 10.36 46.18 10.64 ;
  LAYER M2 ;
        RECT 45.84 9.94 47.04 10.22 ;
  LAYER M2 ;
        RECT 45.41 13.72 47.47 14 ;
  LAYER M1 ;
        RECT 37.715 11.255 37.965 14.785 ;
  LAYER M1 ;
        RECT 37.715 9.995 37.965 11.005 ;
  LAYER M1 ;
        RECT 37.715 7.895 37.965 8.905 ;
  LAYER M1 ;
        RECT 43.735 11.255 43.985 14.785 ;
  LAYER M1 ;
        RECT 31.695 11.255 31.945 14.785 ;
  LAYER M2 ;
        RECT 31.65 14.56 44.03 14.84 ;
  LAYER M2 ;
        RECT 37.24 8.26 38.44 8.54 ;
  LAYER M2 ;
        RECT 37.24 14.14 38.44 14.42 ;
  LAYER M2 ;
        RECT 37.67 10.36 38.87 10.64 ;
  LAYER M3 ;
        RECT 37.27 8.24 37.55 14.86 ;
  LAYER M1 ;
        RECT 54.915 11.255 55.165 14.785 ;
  LAYER M1 ;
        RECT 54.915 9.995 55.165 11.005 ;
  LAYER M1 ;
        RECT 54.915 7.895 55.165 8.905 ;
  LAYER M1 ;
        RECT 48.895 11.255 49.145 14.785 ;
  LAYER M1 ;
        RECT 60.935 11.255 61.185 14.785 ;
  LAYER M2 ;
        RECT 48.85 14.56 61.23 14.84 ;
  LAYER M2 ;
        RECT 54.44 8.26 55.64 8.54 ;
  LAYER M2 ;
        RECT 54.44 14.14 55.64 14.42 ;
  LAYER M2 ;
        RECT 54.01 10.36 55.21 10.64 ;
  LAYER M3 ;
        RECT 55.33 8.24 55.61 14.86 ;
  LAYER M3 ;
        RECT 45.87 22.94 46.15 27.46 ;
  LAYER M2 ;
        RECT 44.98 19.6 46.18 19.88 ;
  LAYER M2 ;
        RECT 37.67 19.6 38.87 19.88 ;
  LAYER M3 ;
        RECT 45.87 19.74 46.15 23.1 ;
  LAYER M2 ;
        RECT 45.85 19.6 46.17 19.88 ;
  LAYER M2 ;
        RECT 38.7 19.6 45.15 19.88 ;
  LAYER M2 ;
        RECT 45.85 19.6 46.17 19.88 ;
  LAYER M3 ;
        RECT 45.87 19.58 46.15 19.9 ;
  LAYER M2 ;
        RECT 45.85 19.6 46.17 19.88 ;
  LAYER M3 ;
        RECT 45.87 19.58 46.15 19.9 ;
  LAYER M2 ;
        RECT 45.85 19.6 46.17 19.88 ;
  LAYER M3 ;
        RECT 45.87 19.58 46.15 19.9 ;
  LAYER M2 ;
        RECT 45.85 19.6 46.17 19.88 ;
  LAYER M3 ;
        RECT 45.87 19.58 46.15 19.9 ;
  LAYER M3 ;
        RECT 46.3 23.36 46.58 27.88 ;
  LAYER M2 ;
        RECT 45.84 20.02 47.04 20.3 ;
  LAYER M2 ;
        RECT 54.01 19.6 55.21 19.88 ;
  LAYER M3 ;
        RECT 46.3 20.16 46.58 23.52 ;
  LAYER M2 ;
        RECT 46.28 20.02 46.6 20.3 ;
  LAYER M2 ;
        RECT 46.71 20.02 47.03 20.3 ;
  LAYER M3 ;
        RECT 46.73 19.74 47.01 20.16 ;
  LAYER M2 ;
        RECT 46.87 19.6 54.18 19.88 ;
  LAYER M2 ;
        RECT 46.28 20.02 46.6 20.3 ;
  LAYER M3 ;
        RECT 46.3 20 46.58 20.32 ;
  LAYER M2 ;
        RECT 46.28 20.02 46.6 20.3 ;
  LAYER M3 ;
        RECT 46.3 20 46.58 20.32 ;
  LAYER M2 ;
        RECT 46.28 20.02 46.6 20.3 ;
  LAYER M3 ;
        RECT 46.3 20 46.58 20.32 ;
  LAYER M2 ;
        RECT 46.71 19.6 47.03 19.88 ;
  LAYER M3 ;
        RECT 46.73 19.58 47.01 19.9 ;
  LAYER M2 ;
        RECT 46.71 20.02 47.03 20.3 ;
  LAYER M3 ;
        RECT 46.73 20 47.01 20.32 ;
  LAYER M2 ;
        RECT 46.28 20.02 46.6 20.3 ;
  LAYER M3 ;
        RECT 46.3 20 46.58 20.32 ;
  LAYER M2 ;
        RECT 46.71 19.6 47.03 19.88 ;
  LAYER M3 ;
        RECT 46.73 19.58 47.01 19.9 ;
  LAYER M2 ;
        RECT 46.71 20.02 47.03 20.3 ;
  LAYER M3 ;
        RECT 46.73 20 47.01 20.32 ;
  LAYER M1 ;
        RECT 45.885 23.015 46.135 26.545 ;
  LAYER M1 ;
        RECT 45.885 26.795 46.135 27.805 ;
  LAYER M1 ;
        RECT 45.885 28.895 46.135 29.905 ;
  LAYER M1 ;
        RECT 45.455 23.015 45.705 26.545 ;
  LAYER M1 ;
        RECT 46.315 23.015 46.565 26.545 ;
  LAYER M1 ;
        RECT 46.745 23.015 46.995 26.545 ;
  LAYER M1 ;
        RECT 46.745 26.795 46.995 27.805 ;
  LAYER M1 ;
        RECT 46.745 28.895 46.995 29.905 ;
  LAYER M1 ;
        RECT 47.175 23.015 47.425 26.545 ;
  LAYER M2 ;
        RECT 44.98 22.96 46.18 23.24 ;
  LAYER M2 ;
        RECT 45.84 27.16 47.04 27.44 ;
  LAYER M2 ;
        RECT 45.84 23.38 47.04 23.66 ;
  LAYER M2 ;
        RECT 45.41 27.58 46.61 27.86 ;
  LAYER M2 ;
        RECT 45.84 29.26 47.04 29.54 ;
  LAYER M3 ;
        RECT 45.87 22.94 46.15 27.46 ;
  LAYER M3 ;
        RECT 46.3 23.36 46.58 27.88 ;
  LAYER M2 ;
        RECT 45.41 23.8 47.47 24.08 ;
  LAYER M1 ;
        RECT 45.885 15.455 46.135 18.985 ;
  LAYER M1 ;
        RECT 45.885 19.235 46.135 20.245 ;
  LAYER M1 ;
        RECT 45.885 21.335 46.135 22.345 ;
  LAYER M1 ;
        RECT 45.455 15.455 45.705 18.985 ;
  LAYER M1 ;
        RECT 46.315 15.455 46.565 18.985 ;
  LAYER M1 ;
        RECT 46.745 15.455 46.995 18.985 ;
  LAYER M1 ;
        RECT 46.745 19.235 46.995 20.245 ;
  LAYER M1 ;
        RECT 46.745 21.335 46.995 22.345 ;
  LAYER M1 ;
        RECT 47.175 15.455 47.425 18.985 ;
  LAYER M2 ;
        RECT 45.84 21.7 47.04 21.98 ;
  LAYER M2 ;
        RECT 44.98 15.4 46.18 15.68 ;
  LAYER M2 ;
        RECT 45.84 15.82 47.04 16.1 ;
  LAYER M2 ;
        RECT 44.98 19.6 46.18 19.88 ;
  LAYER M2 ;
        RECT 45.84 20.02 47.04 20.3 ;
  LAYER M2 ;
        RECT 45.41 16.24 47.47 16.52 ;
  LAYER M1 ;
        RECT 37.715 15.455 37.965 18.985 ;
  LAYER M1 ;
        RECT 37.715 19.235 37.965 20.245 ;
  LAYER M1 ;
        RECT 37.715 21.335 37.965 22.345 ;
  LAYER M1 ;
        RECT 43.735 15.455 43.985 18.985 ;
  LAYER M1 ;
        RECT 31.695 15.455 31.945 18.985 ;
  LAYER M2 ;
        RECT 31.65 15.4 44.03 15.68 ;
  LAYER M2 ;
        RECT 37.24 21.7 38.44 21.98 ;
  LAYER M2 ;
        RECT 37.24 15.82 38.44 16.1 ;
  LAYER M2 ;
        RECT 37.67 19.6 38.87 19.88 ;
  LAYER M3 ;
        RECT 37.27 15.38 37.55 22 ;
  LAYER M1 ;
        RECT 54.915 15.455 55.165 18.985 ;
  LAYER M1 ;
        RECT 54.915 19.235 55.165 20.245 ;
  LAYER M1 ;
        RECT 54.915 21.335 55.165 22.345 ;
  LAYER M1 ;
        RECT 48.895 15.455 49.145 18.985 ;
  LAYER M1 ;
        RECT 60.935 15.455 61.185 18.985 ;
  LAYER M2 ;
        RECT 48.85 15.4 61.23 15.68 ;
  LAYER M2 ;
        RECT 54.44 21.7 55.64 21.98 ;
  LAYER M2 ;
        RECT 54.44 15.82 55.64 16.1 ;
  LAYER M2 ;
        RECT 54.01 19.6 55.21 19.88 ;
  LAYER M3 ;
        RECT 55.33 15.38 55.61 22 ;
  END 
END DCDC_CONV2TO1_1
