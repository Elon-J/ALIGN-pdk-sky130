MACRO CCP_PMOS_58853955_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CCP_PMOS_58853955_X1_Y1 0 0 ;
  SIZE 3440 BY 7560 ;
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1150 260 1430 4780 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 680 1860 5200 ;
    END
  END DB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2010 1100 2290 6880 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 7225 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M2 ;
      RECT 260 280 1460 560 ;
    LAYER M2 ;
      RECT 1120 4480 2320 4760 ;
    LAYER M2 ;
      RECT 1120 700 2320 980 ;
    LAYER M2 ;
      RECT 690 4900 1890 5180 ;
    LAYER M2 ;
      RECT 1120 6580 2320 6860 ;
    LAYER M2 ;
      RECT 690 1120 2750 1400 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4955 1375 5125 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 2065 755 2235 925 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 1635 1175 1805 1345 ;
    LAYER V1 ;
      RECT 2495 1175 2665 1345 ;
    LAYER V2 ;
      RECT 1215 345 1365 495 ;
    LAYER V2 ;
      RECT 1215 4545 1365 4695 ;
    LAYER V2 ;
      RECT 1645 765 1795 915 ;
    LAYER V2 ;
      RECT 1645 4965 1795 5115 ;
    LAYER V2 ;
      RECT 2075 1185 2225 1335 ;
    LAYER V2 ;
      RECT 2075 6645 2225 6795 ;
    LAYER V0 ;
      RECT 1205 2705 1375 2875 ;
    LAYER V0 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V0 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V0 ;
      RECT 775 2705 945 2875 ;
    LAYER V0 ;
      RECT 1635 2705 1805 2875 ;
    LAYER V0 ;
      RECT 1635 2705 1805 2875 ;
    LAYER V0 ;
      RECT 2065 2705 2235 2875 ;
    LAYER V0 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V0 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V0 ;
      RECT 2495 2705 2665 2875 ;
  END
END CCP_PMOS_58853955_X1_Y1
MACRO CMC_PMOS_23131506_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CMC_PMOS_23131506_X1_Y1 0 0 ;
  SIZE 3440 BY 7560 ;
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260 280 1460 560 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 700 2320 980 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 4480 2320 4760 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2440 1100 2720 6880 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 7225 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M2 ;
      RECT 1120 6580 2750 6860 ;
    LAYER M2 ;
      RECT 690 1120 2750 1400 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 2065 755 2235 925 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 1635 1175 1805 1345 ;
    LAYER V1 ;
      RECT 2495 1175 2665 1345 ;
    LAYER V2 ;
      RECT 2505 1185 2655 1335 ;
    LAYER V2 ;
      RECT 2505 6645 2655 6795 ;
    LAYER V0 ;
      RECT 1205 2705 1375 2875 ;
    LAYER V0 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V0 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V0 ;
      RECT 775 2705 945 2875 ;
    LAYER V0 ;
      RECT 1635 2705 1805 2875 ;
    LAYER V0 ;
      RECT 1635 2705 1805 2875 ;
    LAYER V0 ;
      RECT 2065 2705 2235 2875 ;
    LAYER V0 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V0 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V0 ;
      RECT 2495 2705 2665 2875 ;
  END
END CMC_PMOS_23131506_X1_Y1
MACRO CCP_S_NMOS_B_5782581_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CCP_S_NMOS_B_5782581_X1_Y1 0 0 ;
  SIZE 6020 BY 7560 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 6580 4900 6860 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2870 260 3150 4780 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 3300 680 3580 5200 ;
    END
  END DB
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 690 1120 1890 1400 ;
    END
  END SA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4130 1540 5330 1820 ;
    END
  END SB
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 7225 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M2 ;
      RECT 1120 280 3180 560 ;
    LAYER M2 ;
      RECT 2840 4480 4900 4760 ;
    LAYER M2 ;
      RECT 3270 700 4900 980 ;
    LAYER M2 ;
      RECT 1120 4900 3610 5180 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4955 1375 5125 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 4645 755 4815 925 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6635 4815 6805 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 1635 1175 1805 1345 ;
    LAYER V1 ;
      RECT 4215 1595 4385 1765 ;
    LAYER V1 ;
      RECT 5075 1595 5245 1765 ;
    LAYER V2 ;
      RECT 2935 345 3085 495 ;
    LAYER V2 ;
      RECT 2935 4545 3085 4695 ;
    LAYER V2 ;
      RECT 3365 765 3515 915 ;
    LAYER V2 ;
      RECT 3365 4965 3515 5115 ;
    LAYER V0 ;
      RECT 1205 2705 1375 2875 ;
    LAYER V0 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V0 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V0 ;
      RECT 775 2705 945 2875 ;
    LAYER V0 ;
      RECT 1635 2705 1805 2875 ;
    LAYER V0 ;
      RECT 4645 2705 4815 2875 ;
    LAYER V0 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V0 ;
      RECT 4645 6635 4815 6805 ;
    LAYER V0 ;
      RECT 4215 2705 4385 2875 ;
    LAYER V0 ;
      RECT 5075 2705 5245 2875 ;
  END
END CCP_S_NMOS_B_5782581_X1_Y1
MACRO DP_NMOS_B_93310865_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_B_93310865_X1_Y1 0 0 ;
  SIZE 3440 BY 7560 ;
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 6580 2320 6860 ;
    END
  END B
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260 280 1460 560 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 700 2320 980 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260 4480 1460 4760 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1120 4900 2320 5180 ;
    END
  END GB
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 690 1120 2750 1400 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 7225 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 2065 755 2235 925 ;
    LAYER V1 ;
      RECT 2065 4955 2235 5125 ;
    LAYER V1 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V1 ;
      RECT 775 1175 945 1345 ;
    LAYER V1 ;
      RECT 1635 1175 1805 1345 ;
    LAYER V1 ;
      RECT 2495 1175 2665 1345 ;
    LAYER V0 ;
      RECT 1205 2705 1375 2875 ;
    LAYER V0 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V0 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V0 ;
      RECT 775 2705 945 2875 ;
    LAYER V0 ;
      RECT 1635 2705 1805 2875 ;
    LAYER V0 ;
      RECT 1635 2705 1805 2875 ;
    LAYER V0 ;
      RECT 2065 2705 2235 2875 ;
    LAYER V0 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V0 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V0 ;
      RECT 2495 2705 2665 2875 ;
  END
END DP_NMOS_B_93310865_X1_Y1
MACRO NMOS_S_93862694_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_93862694_X1_Y1 0 0 ;
  SIZE 2580 BY 7560 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260 280 1460 560 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260 4480 1460 4760 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 680 1860 6880 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M2 ;
      RECT 690 6580 1890 6860 ;
    LAYER M2 ;
      RECT 690 700 1890 980 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V2 ;
      RECT 1645 765 1795 915 ;
    LAYER V2 ;
      RECT 1645 6645 1795 6795 ;
    LAYER V0 ;
      RECT 1205 2495 1375 2665 ;
    LAYER V0 ;
      RECT 1205 2835 1375 3005 ;
    LAYER V0 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V0 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V0 ;
      RECT 775 2495 945 2665 ;
    LAYER V0 ;
      RECT 775 2835 945 3005 ;
    LAYER V0 ;
      RECT 1635 2495 1805 2665 ;
    LAYER V0 ;
      RECT 1635 2835 1805 3005 ;
  END
END NMOS_S_93862694_X1_Y1
