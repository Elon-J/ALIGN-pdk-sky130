MACRO DCDC_HUNIT_CONV2TO1
  ORIGIN 0 0 ;
  FOREIGN DCDC_HUNIT_CONV2TO1 0 0 ;
  SIZE 31.82 BY 31.5 ;
  PIN CLK1B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 6.31 8.66 6.59 15.28 ;
    END
  END CLK1B
  PIN CLK0B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 25.23 8.66 25.51 15.28 ;
    END
  END CLK0B
  PIN VHIGH
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.88 6.16 16.94 6.44 ;
      LAYER M2 ;
        RECT 14.88 14.14 16.94 14.42 ;
      LAYER M2 ;
        RECT 14.89 6.16 15.21 6.44 ;
      LAYER M3 ;
        RECT 14.91 6.3 15.19 14.28 ;
      LAYER M2 ;
        RECT 14.89 14.14 15.21 14.42 ;
    END
  END VHIGH
  PIN Y0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 16.17 14.98 17.37 15.26 ;
      LAYER M2 ;
        RECT 16.17 16.24 17.37 16.52 ;
      LAYER M2 ;
        RECT 16.61 14.98 16.93 15.26 ;
      LAYER M3 ;
        RECT 16.63 15.12 16.91 16.38 ;
      LAYER M2 ;
        RECT 16.61 16.24 16.93 16.52 ;
    END
  END Y0
  PIN Y1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.31 14.56 16.51 14.84 ;
      LAYER M2 ;
        RECT 15.31 16.66 16.51 16.94 ;
      LAYER M2 ;
        RECT 15.75 14.56 16.07 14.84 ;
      LAYER M3 ;
        RECT 15.77 14.7 16.05 16.8 ;
      LAYER M2 ;
        RECT 15.75 16.66 16.07 16.94 ;
    END
  END Y1
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.31 0.7 16.51 0.98 ;
      LAYER M2 ;
        RECT 15.31 8.68 16.51 8.96 ;
      LAYER M2 ;
        RECT 15.32 0.7 15.64 0.98 ;
      LAYER M3 ;
        RECT 15.34 0.84 15.62 8.82 ;
      LAYER M2 ;
        RECT 15.32 8.68 15.64 8.96 ;
    END
  END VPWR
  PIN CLK0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 6.31 16.22 6.59 22.84 ;
    END
  END CLK0
  PIN CLK1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 25.23 16.22 25.51 22.84 ;
    END
  END CLK1
  PIN VLOW
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.88 25.06 16.94 25.34 ;
      LAYER M2 ;
        RECT 14.88 17.08 16.94 17.36 ;
      LAYER M2 ;
        RECT 14.89 25.06 15.21 25.34 ;
      LAYER M3 ;
        RECT 14.91 17.22 15.19 25.2 ;
      LAYER M2 ;
        RECT 14.89 17.08 15.21 17.36 ;
    END
  END VLOW
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.31 30.52 16.51 30.8 ;
      LAYER M2 ;
        RECT 15.31 22.54 16.51 22.82 ;
      LAYER M2 ;
        RECT 15.32 30.52 15.64 30.8 ;
      LAYER M3 ;
        RECT 15.34 22.68 15.62 30.66 ;
      LAYER M2 ;
        RECT 15.32 22.54 15.64 22.82 ;
    END
  END VGND
  OBS 
  LAYER M3 ;
        RECT 16.2 2.78 16.48 7.3 ;
  LAYER M2 ;
        RECT 16.17 10.78 17.37 11.06 ;
  LAYER M2 ;
        RECT 23.91 10.78 25.11 11.06 ;
  LAYER M3 ;
        RECT 16.2 7.14 16.48 10.92 ;
  LAYER M2 ;
        RECT 16.18 10.78 16.5 11.06 ;
  LAYER M2 ;
        RECT 17.2 10.78 24.08 11.06 ;
  LAYER M2 ;
        RECT 16.18 10.78 16.5 11.06 ;
  LAYER M3 ;
        RECT 16.2 10.76 16.48 11.08 ;
  LAYER M2 ;
        RECT 16.18 10.78 16.5 11.06 ;
  LAYER M3 ;
        RECT 16.2 10.76 16.48 11.08 ;
  LAYER M2 ;
        RECT 16.18 10.78 16.5 11.06 ;
  LAYER M3 ;
        RECT 16.2 10.76 16.48 11.08 ;
  LAYER M2 ;
        RECT 16.18 10.78 16.5 11.06 ;
  LAYER M3 ;
        RECT 16.2 10.76 16.48 11.08 ;
  LAYER M3 ;
        RECT 15.77 2.36 16.05 6.88 ;
  LAYER M2 ;
        RECT 15.31 10.36 16.51 10.64 ;
  LAYER M2 ;
        RECT 6.71 10.78 7.91 11.06 ;
  LAYER M3 ;
        RECT 15.77 6.72 16.05 10.5 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M2 ;
        RECT 15.32 10.36 15.64 10.64 ;
  LAYER M3 ;
        RECT 15.34 10.5 15.62 10.92 ;
  LAYER M2 ;
        RECT 7.74 10.78 15.48 11.06 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M2 ;
        RECT 15.32 10.36 15.64 10.64 ;
  LAYER M3 ;
        RECT 15.34 10.34 15.62 10.66 ;
  LAYER M2 ;
        RECT 15.32 10.78 15.64 11.06 ;
  LAYER M3 ;
        RECT 15.34 10.76 15.62 11.08 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M2 ;
        RECT 15.32 10.36 15.64 10.64 ;
  LAYER M3 ;
        RECT 15.34 10.34 15.62 10.66 ;
  LAYER M2 ;
        RECT 15.32 10.78 15.64 11.06 ;
  LAYER M3 ;
        RECT 15.34 10.76 15.62 11.08 ;
  LAYER M2 ;
        RECT 15.75 10.36 16.07 10.64 ;
  LAYER M3 ;
        RECT 15.77 10.34 16.05 10.66 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 16.215 2.435 16.465 3.445 ;
  LAYER M1 ;
        RECT 16.215 0.335 16.465 1.345 ;
  LAYER M1 ;
        RECT 16.645 3.695 16.895 7.225 ;
  LAYER M1 ;
        RECT 15.785 3.695 16.035 7.225 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M1 ;
        RECT 15.355 2.435 15.605 3.445 ;
  LAYER M1 ;
        RECT 15.355 0.335 15.605 1.345 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M2 ;
        RECT 16.17 7 17.37 7.28 ;
  LAYER M2 ;
        RECT 15.31 2.8 16.51 3.08 ;
  LAYER M2 ;
        RECT 15.31 6.58 16.51 6.86 ;
  LAYER M2 ;
        RECT 15.74 2.38 16.94 2.66 ;
  LAYER M2 ;
        RECT 15.31 0.7 16.51 0.98 ;
  LAYER M3 ;
        RECT 16.2 2.78 16.48 7.3 ;
  LAYER M3 ;
        RECT 15.77 2.36 16.05 6.88 ;
  LAYER M2 ;
        RECT 14.88 6.16 16.94 6.44 ;
  LAYER M1 ;
        RECT 16.215 11.675 16.465 15.205 ;
  LAYER M1 ;
        RECT 16.215 10.415 16.465 11.425 ;
  LAYER M1 ;
        RECT 16.215 8.315 16.465 9.325 ;
  LAYER M1 ;
        RECT 16.645 11.675 16.895 15.205 ;
  LAYER M1 ;
        RECT 15.785 11.675 16.035 15.205 ;
  LAYER M1 ;
        RECT 15.355 11.675 15.605 15.205 ;
  LAYER M1 ;
        RECT 15.355 10.415 15.605 11.425 ;
  LAYER M1 ;
        RECT 15.355 8.315 15.605 9.325 ;
  LAYER M1 ;
        RECT 14.925 11.675 15.175 15.205 ;
  LAYER M2 ;
        RECT 15.31 8.68 16.51 8.96 ;
  LAYER M2 ;
        RECT 16.17 14.98 17.37 15.26 ;
  LAYER M2 ;
        RECT 15.31 14.56 16.51 14.84 ;
  LAYER M2 ;
        RECT 16.17 10.78 17.37 11.06 ;
  LAYER M2 ;
        RECT 15.31 10.36 16.51 10.64 ;
  LAYER M2 ;
        RECT 14.88 14.14 16.94 14.42 ;
  LAYER M1 ;
        RECT 24.815 11.675 25.065 15.205 ;
  LAYER M1 ;
        RECT 24.815 10.415 25.065 11.425 ;
  LAYER M1 ;
        RECT 24.815 8.315 25.065 9.325 ;
  LAYER M1 ;
        RECT 18.795 11.675 19.045 15.205 ;
  LAYER M1 ;
        RECT 30.835 11.675 31.085 15.205 ;
  LAYER M2 ;
        RECT 24.34 14.98 25.54 15.26 ;
  LAYER M2 ;
        RECT 18.75 14.56 31.13 14.84 ;
  LAYER M2 ;
        RECT 24.34 8.68 25.54 8.96 ;
  LAYER M2 ;
        RECT 23.91 10.78 25.11 11.06 ;
  LAYER M3 ;
        RECT 25.23 8.66 25.51 15.28 ;
  LAYER M1 ;
        RECT 6.755 11.675 7.005 15.205 ;
  LAYER M1 ;
        RECT 6.755 10.415 7.005 11.425 ;
  LAYER M1 ;
        RECT 6.755 8.315 7.005 9.325 ;
  LAYER M1 ;
        RECT 12.775 11.675 13.025 15.205 ;
  LAYER M1 ;
        RECT 0.735 11.675 0.985 15.205 ;
  LAYER M2 ;
        RECT 6.28 14.98 7.48 15.26 ;
  LAYER M2 ;
        RECT 0.69 14.56 13.07 14.84 ;
  LAYER M2 ;
        RECT 6.28 8.68 7.48 8.96 ;
  LAYER M2 ;
        RECT 6.71 10.78 7.91 11.06 ;
  LAYER M3 ;
        RECT 6.31 8.66 6.59 15.28 ;
  LAYER M3 ;
        RECT 16.2 24.2 16.48 28.72 ;
  LAYER M2 ;
        RECT 16.17 20.44 17.37 20.72 ;
  LAYER M2 ;
        RECT 23.91 20.44 25.11 20.72 ;
  LAYER M3 ;
        RECT 16.2 20.58 16.48 24.36 ;
  LAYER M2 ;
        RECT 16.18 20.44 16.5 20.72 ;
  LAYER M2 ;
        RECT 17.2 20.44 24.08 20.72 ;
  LAYER M2 ;
        RECT 16.18 20.44 16.5 20.72 ;
  LAYER M3 ;
        RECT 16.2 20.42 16.48 20.74 ;
  LAYER M2 ;
        RECT 16.18 20.44 16.5 20.72 ;
  LAYER M3 ;
        RECT 16.2 20.42 16.48 20.74 ;
  LAYER M2 ;
        RECT 16.18 20.44 16.5 20.72 ;
  LAYER M3 ;
        RECT 16.2 20.42 16.48 20.74 ;
  LAYER M2 ;
        RECT 16.18 20.44 16.5 20.72 ;
  LAYER M3 ;
        RECT 16.2 20.42 16.48 20.74 ;
  LAYER M3 ;
        RECT 15.77 24.62 16.05 29.14 ;
  LAYER M2 ;
        RECT 15.31 20.86 16.51 21.14 ;
  LAYER M2 ;
        RECT 6.71 20.44 7.91 20.72 ;
  LAYER M3 ;
        RECT 15.77 21 16.05 24.78 ;
  LAYER M2 ;
        RECT 15.75 20.86 16.07 21.14 ;
  LAYER M2 ;
        RECT 15.32 20.86 15.64 21.14 ;
  LAYER M3 ;
        RECT 15.34 20.58 15.62 21 ;
  LAYER M2 ;
        RECT 7.74 20.44 15.48 20.72 ;
  LAYER M2 ;
        RECT 15.75 20.86 16.07 21.14 ;
  LAYER M3 ;
        RECT 15.77 20.84 16.05 21.16 ;
  LAYER M2 ;
        RECT 15.75 20.86 16.07 21.14 ;
  LAYER M3 ;
        RECT 15.77 20.84 16.05 21.16 ;
  LAYER M2 ;
        RECT 15.32 20.86 15.64 21.14 ;
  LAYER M3 ;
        RECT 15.34 20.84 15.62 21.16 ;
  LAYER M2 ;
        RECT 15.32 20.44 15.64 20.72 ;
  LAYER M3 ;
        RECT 15.34 20.42 15.62 20.74 ;
  LAYER M2 ;
        RECT 15.75 20.86 16.07 21.14 ;
  LAYER M3 ;
        RECT 15.77 20.84 16.05 21.16 ;
  LAYER M2 ;
        RECT 15.32 20.86 15.64 21.14 ;
  LAYER M3 ;
        RECT 15.34 20.84 15.62 21.16 ;
  LAYER M2 ;
        RECT 15.32 20.44 15.64 20.72 ;
  LAYER M3 ;
        RECT 15.34 20.42 15.62 20.74 ;
  LAYER M2 ;
        RECT 15.75 20.86 16.07 21.14 ;
  LAYER M3 ;
        RECT 15.77 20.84 16.05 21.16 ;
  LAYER M1 ;
        RECT 16.215 24.275 16.465 27.805 ;
  LAYER M1 ;
        RECT 16.215 28.055 16.465 29.065 ;
  LAYER M1 ;
        RECT 16.215 30.155 16.465 31.165 ;
  LAYER M1 ;
        RECT 16.645 24.275 16.895 27.805 ;
  LAYER M1 ;
        RECT 15.785 24.275 16.035 27.805 ;
  LAYER M1 ;
        RECT 15.355 24.275 15.605 27.805 ;
  LAYER M1 ;
        RECT 15.355 28.055 15.605 29.065 ;
  LAYER M1 ;
        RECT 15.355 30.155 15.605 31.165 ;
  LAYER M1 ;
        RECT 14.925 24.275 15.175 27.805 ;
  LAYER M2 ;
        RECT 16.17 24.22 17.37 24.5 ;
  LAYER M2 ;
        RECT 15.31 28.42 16.51 28.7 ;
  LAYER M2 ;
        RECT 15.31 24.64 16.51 24.92 ;
  LAYER M2 ;
        RECT 15.74 28.84 16.94 29.12 ;
  LAYER M2 ;
        RECT 15.31 30.52 16.51 30.8 ;
  LAYER M3 ;
        RECT 16.2 24.2 16.48 28.72 ;
  LAYER M3 ;
        RECT 15.77 24.62 16.05 29.14 ;
  LAYER M2 ;
        RECT 14.88 25.06 16.94 25.34 ;
  LAYER M1 ;
        RECT 16.215 16.295 16.465 19.825 ;
  LAYER M1 ;
        RECT 16.215 20.075 16.465 21.085 ;
  LAYER M1 ;
        RECT 16.215 22.175 16.465 23.185 ;
  LAYER M1 ;
        RECT 16.645 16.295 16.895 19.825 ;
  LAYER M1 ;
        RECT 15.785 16.295 16.035 19.825 ;
  LAYER M1 ;
        RECT 15.355 16.295 15.605 19.825 ;
  LAYER M1 ;
        RECT 15.355 20.075 15.605 21.085 ;
  LAYER M1 ;
        RECT 15.355 22.175 15.605 23.185 ;
  LAYER M1 ;
        RECT 14.925 16.295 15.175 19.825 ;
  LAYER M2 ;
        RECT 15.31 22.54 16.51 22.82 ;
  LAYER M2 ;
        RECT 16.17 16.24 17.37 16.52 ;
  LAYER M2 ;
        RECT 15.31 16.66 16.51 16.94 ;
  LAYER M2 ;
        RECT 16.17 20.44 17.37 20.72 ;
  LAYER M2 ;
        RECT 15.31 20.86 16.51 21.14 ;
  LAYER M2 ;
        RECT 14.88 17.08 16.94 17.36 ;
  LAYER M1 ;
        RECT 24.815 16.295 25.065 19.825 ;
  LAYER M1 ;
        RECT 24.815 20.075 25.065 21.085 ;
  LAYER M1 ;
        RECT 24.815 22.175 25.065 23.185 ;
  LAYER M1 ;
        RECT 18.795 16.295 19.045 19.825 ;
  LAYER M1 ;
        RECT 30.835 16.295 31.085 19.825 ;
  LAYER M2 ;
        RECT 24.34 16.24 25.54 16.52 ;
  LAYER M2 ;
        RECT 18.75 16.66 31.13 16.94 ;
  LAYER M2 ;
        RECT 24.34 22.54 25.54 22.82 ;
  LAYER M2 ;
        RECT 23.91 20.44 25.11 20.72 ;
  LAYER M3 ;
        RECT 25.23 16.22 25.51 22.84 ;
  LAYER M1 ;
        RECT 6.755 16.295 7.005 19.825 ;
  LAYER M1 ;
        RECT 6.755 20.075 7.005 21.085 ;
  LAYER M1 ;
        RECT 6.755 22.175 7.005 23.185 ;
  LAYER M1 ;
        RECT 12.775 16.295 13.025 19.825 ;
  LAYER M1 ;
        RECT 0.735 16.295 0.985 19.825 ;
  LAYER M2 ;
        RECT 6.28 16.24 7.48 16.52 ;
  LAYER M2 ;
        RECT 0.69 16.66 13.07 16.94 ;
  LAYER M2 ;
        RECT 6.28 22.54 7.48 22.82 ;
  LAYER M2 ;
        RECT 6.71 20.44 7.91 20.72 ;
  LAYER M3 ;
        RECT 6.31 16.22 6.59 22.84 ;
  END 
END DCDC_HUNIT_CONV2TO1
