MACRO DCDC_XSW_PMOS
  ORIGIN 0 0 ;
  FOREIGN DCDC_XSW_PMOS 0 0 ;
  SIZE 30.96 BY 15.12 ;
  PIN VPB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.88 14.14 16.08 14.42 ;
      LAYER M2 ;
        RECT 14.88 6.58 16.08 6.86 ;
      LAYER M2 ;
        RECT 14.89 14.14 15.21 14.42 ;
      LAYER M3 ;
        RECT 14.91 6.72 15.19 14.28 ;
      LAYER M2 ;
        RECT 14.89 6.58 15.21 6.86 ;
    END
  END VPB
  PIN VIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.45 8.68 16.51 8.96 ;
      LAYER M2 ;
        RECT 14.45 1.12 16.51 1.4 ;
      LAYER M2 ;
        RECT 14.46 8.68 14.78 8.96 ;
      LAYER M3 ;
        RECT 14.48 1.26 14.76 8.82 ;
      LAYER M2 ;
        RECT 14.46 1.12 14.78 1.4 ;
    END
  END VIN
  PIN VOUT0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.74 0.28 16.94 0.56 ;
    END
  END VOUT0
  PIN VOUT1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.88 0.7 16.08 0.98 ;
    END
  END VOUT1
  PIN CLKB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 24.37 0.26 24.65 6.88 ;
    END
  END CLKB
  PIN CLK
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 6.31 0.26 6.59 6.88 ;
    END
  END CLK
  OBS 
  LAYER M3 ;
        RECT 15.77 7.82 16.05 12.34 ;
  LAYER M2 ;
        RECT 15.74 4.48 16.94 4.76 ;
  LAYER M2 ;
        RECT 23.05 4.48 24.25 4.76 ;
  LAYER M3 ;
        RECT 15.77 4.62 16.05 7.98 ;
  LAYER M2 ;
        RECT 15.75 4.48 16.07 4.76 ;
  LAYER M2 ;
        RECT 16.77 4.48 23.22 4.76 ;
  LAYER M2 ;
        RECT 15.75 4.48 16.07 4.76 ;
  LAYER M3 ;
        RECT 15.77 4.46 16.05 4.78 ;
  LAYER M2 ;
        RECT 15.75 4.48 16.07 4.76 ;
  LAYER M3 ;
        RECT 15.77 4.46 16.05 4.78 ;
  LAYER M2 ;
        RECT 15.75 4.48 16.07 4.76 ;
  LAYER M3 ;
        RECT 15.77 4.46 16.05 4.78 ;
  LAYER M2 ;
        RECT 15.75 4.48 16.07 4.76 ;
  LAYER M3 ;
        RECT 15.77 4.46 16.05 4.78 ;
  LAYER M3 ;
        RECT 15.34 8.24 15.62 12.76 ;
  LAYER M2 ;
        RECT 14.88 4.9 16.08 5.18 ;
  LAYER M2 ;
        RECT 6.71 4.48 7.91 4.76 ;
  LAYER M3 ;
        RECT 15.34 5.04 15.62 8.4 ;
  LAYER M2 ;
        RECT 15.32 4.9 15.64 5.18 ;
  LAYER M2 ;
        RECT 14.89 4.9 15.21 5.18 ;
  LAYER M3 ;
        RECT 14.91 4.62 15.19 5.04 ;
  LAYER M2 ;
        RECT 7.74 4.48 15.05 4.76 ;
  LAYER M2 ;
        RECT 15.32 4.9 15.64 5.18 ;
  LAYER M3 ;
        RECT 15.34 4.88 15.62 5.2 ;
  LAYER M2 ;
        RECT 15.32 4.9 15.64 5.18 ;
  LAYER M3 ;
        RECT 15.34 4.88 15.62 5.2 ;
  LAYER M2 ;
        RECT 14.89 4.9 15.21 5.18 ;
  LAYER M3 ;
        RECT 14.91 4.88 15.19 5.2 ;
  LAYER M2 ;
        RECT 14.89 4.48 15.21 4.76 ;
  LAYER M3 ;
        RECT 14.91 4.46 15.19 4.78 ;
  LAYER M2 ;
        RECT 15.32 4.9 15.64 5.18 ;
  LAYER M3 ;
        RECT 15.34 4.88 15.62 5.2 ;
  LAYER M2 ;
        RECT 14.89 4.9 15.21 5.18 ;
  LAYER M3 ;
        RECT 14.91 4.88 15.19 5.2 ;
  LAYER M2 ;
        RECT 14.89 4.48 15.21 4.76 ;
  LAYER M3 ;
        RECT 14.91 4.46 15.19 4.78 ;
  LAYER M2 ;
        RECT 15.32 4.9 15.64 5.18 ;
  LAYER M3 ;
        RECT 15.34 4.88 15.62 5.2 ;
  LAYER M1 ;
        RECT 15.785 7.895 16.035 11.425 ;
  LAYER M1 ;
        RECT 15.785 11.675 16.035 12.685 ;
  LAYER M1 ;
        RECT 15.785 13.775 16.035 14.785 ;
  LAYER M1 ;
        RECT 16.215 7.895 16.465 11.425 ;
  LAYER M1 ;
        RECT 15.355 7.895 15.605 11.425 ;
  LAYER M1 ;
        RECT 14.925 7.895 15.175 11.425 ;
  LAYER M1 ;
        RECT 14.925 11.675 15.175 12.685 ;
  LAYER M1 ;
        RECT 14.925 13.775 15.175 14.785 ;
  LAYER M1 ;
        RECT 14.495 7.895 14.745 11.425 ;
  LAYER M2 ;
        RECT 15.74 7.84 16.94 8.12 ;
  LAYER M2 ;
        RECT 14.88 12.04 16.08 12.32 ;
  LAYER M2 ;
        RECT 14.88 8.26 16.08 8.54 ;
  LAYER M2 ;
        RECT 15.31 12.46 16.51 12.74 ;
  LAYER M2 ;
        RECT 14.88 14.14 16.08 14.42 ;
  LAYER M3 ;
        RECT 15.77 7.82 16.05 12.34 ;
  LAYER M3 ;
        RECT 15.34 8.24 15.62 12.76 ;
  LAYER M2 ;
        RECT 14.45 8.68 16.51 8.96 ;
  LAYER M1 ;
        RECT 15.785 0.335 16.035 3.865 ;
  LAYER M1 ;
        RECT 15.785 4.115 16.035 5.125 ;
  LAYER M1 ;
        RECT 15.785 6.215 16.035 7.225 ;
  LAYER M1 ;
        RECT 16.215 0.335 16.465 3.865 ;
  LAYER M1 ;
        RECT 15.355 0.335 15.605 3.865 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 3.865 ;
  LAYER M1 ;
        RECT 14.925 4.115 15.175 5.125 ;
  LAYER M1 ;
        RECT 14.925 6.215 15.175 7.225 ;
  LAYER M1 ;
        RECT 14.495 0.335 14.745 3.865 ;
  LAYER M2 ;
        RECT 14.88 6.58 16.08 6.86 ;
  LAYER M2 ;
        RECT 15.74 0.28 16.94 0.56 ;
  LAYER M2 ;
        RECT 14.88 0.7 16.08 0.98 ;
  LAYER M2 ;
        RECT 15.74 4.48 16.94 4.76 ;
  LAYER M2 ;
        RECT 14.88 4.9 16.08 5.18 ;
  LAYER M2 ;
        RECT 14.45 1.12 16.51 1.4 ;
  LAYER M1 ;
        RECT 23.955 0.335 24.205 3.865 ;
  LAYER M1 ;
        RECT 23.955 4.115 24.205 5.125 ;
  LAYER M1 ;
        RECT 23.955 6.215 24.205 7.225 ;
  LAYER M1 ;
        RECT 17.935 0.335 18.185 3.865 ;
  LAYER M1 ;
        RECT 29.975 0.335 30.225 3.865 ;
  LAYER M2 ;
        RECT 17.89 0.28 30.27 0.56 ;
  LAYER M2 ;
        RECT 23.48 6.58 24.68 6.86 ;
  LAYER M2 ;
        RECT 23.48 0.7 24.68 0.98 ;
  LAYER M2 ;
        RECT 23.05 4.48 24.25 4.76 ;
  LAYER M3 ;
        RECT 24.37 0.26 24.65 6.88 ;
  LAYER M1 ;
        RECT 6.755 0.335 7.005 3.865 ;
  LAYER M1 ;
        RECT 6.755 4.115 7.005 5.125 ;
  LAYER M1 ;
        RECT 6.755 6.215 7.005 7.225 ;
  LAYER M1 ;
        RECT 12.775 0.335 13.025 3.865 ;
  LAYER M1 ;
        RECT 0.735 0.335 0.985 3.865 ;
  LAYER M2 ;
        RECT 0.69 0.28 13.07 0.56 ;
  LAYER M2 ;
        RECT 6.28 6.58 7.48 6.86 ;
  LAYER M2 ;
        RECT 6.28 0.7 7.48 0.98 ;
  LAYER M2 ;
        RECT 6.71 4.48 7.91 4.76 ;
  LAYER M3 ;
        RECT 6.31 0.26 6.59 6.88 ;
  END 
END DCDC_XSW_PMOS
