MACRO CAP_2T_42108783
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN CAP_2T_42108783 0 0 ;
  SIZE 1000001980 BY 16000005420 ;
  PIN MINUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 265 860 1000001285 1660 ;
    END
  END MINUS
  PIN PLUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 265 16000003760 1000001285 16000004560 ;
    END
  END PLUS
  OBS
    LAYER M4 ;
      RECT 860 2370 1000001160 16000002670 ;
    LAYER M4 ;
      RECT 1000000710 16000001440 1000001160 16000003960 ;
    LAYER M5 ;
      RECT 1085 830 1535 3350 ;
    LAYER V4 ;
      RECT 1210 1160 1410 1360 ;
  END
END CAP_2T_42108783
